<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-61.7833,42.7185,228.35,-100.689</PageViewport>
<gate>
<ID>2</ID>
<type>AE_DFF_LOW</type>
<position>43,-44</position>
<input>
<ID>IN_0</ID>4 </input>
<output>
<ID>OUT_0</ID>19 </output>
<input>
<ID>clock</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4</ID>
<type>AE_DFF_LOW</type>
<position>70.5,-45</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>20 </output>
<input>
<ID>clock</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_DFF_LOW</type>
<position>94,-45.5</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>21 </output>
<input>
<ID>clock</ID>3 </input>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8</ID>
<type>AE_DFF_LOW</type>
<position>117.5,-45.5</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>23 </output>
<input>
<ID>clock</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>12,-15</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>12</ID>
<type>BB_CLOCK</type>
<position>26.5,-55</position>
<output>
<ID>CLK</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_INVERTER</type>
<position>25,-1.5</position>
<input>
<ID>IN_0</ID>17 </input>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_AND2</type>
<position>30.5,-18</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_AND2</type>
<position>37.5,-18</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AE_OR2</type>
<position>34,-30</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_AND2</type>
<position>57.5,-18</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_AND2</type>
<position>64.5,-18</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>AE_OR2</type>
<position>61,-30</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_AND2</type>
<position>80,-18</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_AND2</type>
<position>87,-18</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>34</ID>
<type>AE_OR2</type>
<position>83.5,-30</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>GA_LED</type>
<position>49.5,-60</position>
<input>
<ID>N_in3</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>GA_LED</type>
<position>75,-59.5</position>
<input>
<ID>N_in3</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>GA_LED</type>
<position>100,-60</position>
<input>
<ID>N_in3</ID>21 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>GA_LED</type>
<position>122.5,-61</position>
<input>
<ID>N_in3</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_AND2</type>
<position>107,-18.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND2</type>
<position>114,-18.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>AE_OR2</type>
<position>110.5,-30.5</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_TOGGLE</type>
<position>17,-7.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_TOGGLE</type>
<position>130,-14.5</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_LABEL</type>
<position>82.5,22</position>
<gparam>LABEL_TEXT 4-bit PISO (Right/Left')</gparam>
<gparam>TEXT_HEIGHT 6</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>0.5,-14.5</position>
<gparam>LABEL_TEXT Shift Right</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>141.5,-14</position>
<gparam>LABEL_TEXT Shift Left</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14,-15,29.5,-15</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-55,112,-46.5</points>
<intersection>-55 2</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-46.5,114.5,-46.5</points>
<connection>
<GID>8</GID>
<name>clock</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-55,112,-55</points>
<connection>
<GID>12</GID>
<name>CLK</name></connection>
<intersection>40 5</intersection>
<intersection>67.5 4</intersection>
<intersection>91 3</intersection>
<intersection>112 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>91,-55,91,-46.5</points>
<connection>
<GID>6</GID>
<name>clock</name></connection>
<intersection>-55 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>67.5,-55,67.5,-46</points>
<connection>
<GID>4</GID>
<name>clock</name></connection>
<intersection>-55 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>40,-55,40,-45</points>
<connection>
<GID>2</GID>
<name>clock</name></connection>
<intersection>-55 2</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-42,34,-33</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-42,40,-42</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-43,61,-33</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-43,67.5,-43</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-43.5,83.5,-33</points>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-43.5,91,-43.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-43.5,110.5,-33.5</points>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110.5,-43.5,114.5,-43.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>110.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-27,35,-24</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>-24 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>37.5,-24,37.5,-21</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>35,-24,37.5,-24</points>
<intersection>35 0</intersection>
<intersection>37.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-27,33,-24</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>-24 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>30.5,-24,30.5,-21</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-24,33,-24</points>
<intersection>30.5 1</intersection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-27,62,-24</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>-24 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>64.5,-24,64.5,-21</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>62,-24,64.5,-24</points>
<intersection>62 0</intersection>
<intersection>64.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-27,60,-24</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>-24 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>57.5,-24,57.5,-21</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-24,60,-24</points>
<intersection>57.5 1</intersection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-27,84.5,-24</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>-24 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>87,-24,87,-21</points>
<connection>
<GID>33</GID>
<name>OUT</name></connection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-24,87,-24</points>
<intersection>84.5 0</intersection>
<intersection>87 1</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-27,82.5,-24</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<intersection>-24 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>80,-24,80,-21</points>
<connection>
<GID>32</GID>
<name>OUT</name></connection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>80,-24,82.5,-24</points>
<intersection>80 1</intersection>
<intersection>82.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-27.5,109.5,-24.5</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>-24.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>107,-24.5,107,-21.5</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>107,-24.5,109.5,-24.5</points>
<intersection>107 1</intersection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-27.5,111.5,-24.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>-24.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>114,-24.5,114,-21.5</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>111.5,-24.5,114,-24.5</points>
<intersection>111.5 0</intersection>
<intersection>114 1</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-15.5,108,-7.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-7.5,108,-7.5</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<intersection>22 2</intersection>
<intersection>31.5 3</intersection>
<intersection>58.5 4</intersection>
<intersection>81 5</intersection>
<intersection>108 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>22,-7.5,22,-1.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>-7.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>31.5,-15,31.5,-7.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-7.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>58.5,-15,58.5,-7.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>-7.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>81,-15,81,-7.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>-7.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,-15.5,113,-1.5</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-1.5,113,-1.5</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>36.5 2</intersection>
<intersection>63.5 4</intersection>
<intersection>86 3</intersection>
<intersection>113 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>36.5,-15,36.5,-1.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>-1.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>86,-15,86,-1.5</points>
<connection>
<GID>33</GID>
<name>IN_1</name></connection>
<intersection>-1.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>63.5,-15,63.5,-1.5</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>-1.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-42,53,-15</points>
<intersection>-42 1</intersection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-42,53,-42</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>49.5 3</intersection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,-15,56.5,-15</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>53 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>49.5,-59,49.5,-42</points>
<connection>
<GID>36</GID>
<name>N_in3</name></connection>
<intersection>-42 1</intersection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-43,77,10</points>
<intersection>-43 1</intersection>
<intersection>-15 2</intersection>
<intersection>10 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-43,77,-43</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>75 6</intersection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-15,79,-15</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>38.5,10,77,10</points>
<intersection>38.5 5</intersection>
<intersection>77 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>38.5,-15,38.5,10</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>10 4</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>75,-58.5,75,-43</points>
<connection>
<GID>38</GID>
<name>N_in3</name></connection>
<intersection>-43 1</intersection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-43.5,103,5</points>
<intersection>-43.5 1</intersection>
<intersection>-15.5 2</intersection>
<intersection>5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97,-43.5,103,-43.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>100 5</intersection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-15.5,106,-15.5</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>65.5,5,103,5</points>
<intersection>65.5 4</intersection>
<intersection>103 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>65.5,-15,65.5,5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>5 3</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>100,-59,100,-43.5</points>
<connection>
<GID>40</GID>
<name>N_in3</name></connection>
<intersection>-43.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-15.5,115,-14.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-14.5,128,-14.5</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-43.5,124.5,2.5</points>
<intersection>-43.5 4</intersection>
<intersection>2.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>88,2.5,124.5,2.5</points>
<intersection>88 3</intersection>
<intersection>124.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>88,-15,88,2.5</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>2.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>120.5,-43.5,124.5,-43.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>122.5 11</intersection>
<intersection>124.5 0</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>122.5,-60,122.5,-43.5</points>
<connection>
<GID>42</GID>
<name>N_in3</name></connection>
<intersection>-43.5 4</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>-116.6,44.4889,101,-63.0667</PageViewport>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>-2.5,12</position>
<gparam>LABEL_TEXT Universal Shift Resistor</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AE_MUX_4x1</type>
<position>-41,-34.5</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_2</ID>37 </input>
<input>
<ID>IN_3</ID>24 </input>
<input>
<ID>SEL_0</ID>43 </input>
<input>
<ID>SEL_1</ID>42 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>59</ID>
<type>AE_MUX_4x1</type>
<position>-17,-35</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>48 </input>
<input>
<ID>IN_2</ID>38 </input>
<input>
<ID>IN_3</ID>25 </input>
<input>
<ID>SEL_0</ID>43 </input>
<input>
<ID>SEL_1</ID>42 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>60</ID>
<type>AE_MUX_4x1</type>
<position>6,-35.5</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>51 </input>
<input>
<ID>IN_2</ID>39 </input>
<input>
<ID>IN_3</ID>26 </input>
<input>
<ID>SEL_0</ID>43 </input>
<input>
<ID>SEL_1</ID>42 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>61</ID>
<type>AE_MUX_4x1</type>
<position>28.5,-36</position>
<input>
<ID>IN_1</ID>50 </input>
<input>
<ID>IN_2</ID>40 </input>
<input>
<ID>IN_3</ID>27 </input>
<input>
<ID>SEL_0</ID>43 </input>
<input>
<ID>SEL_1</ID>42 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_TOGGLE</type>
<position>-44,-47.5</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_TOGGLE</type>
<position>-20,-47.5</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_TOGGLE</type>
<position>3,-48</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_TOGGLE</type>
<position>25.5,-48</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>77</ID>
<type>BB_CLOCK</type>
<position>-52.5,-22.5</position>
<output>
<ID>CLK</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>79</ID>
<type>AE_DFF_LOW</type>
<position>-36,-11</position>
<output>
<ID>OUTINV_0</ID>48 </output>
<output>
<ID>OUT_0</ID>37 </output>
<input>
<ID>clock</ID>36 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>80</ID>
<type>AE_DFF_LOW</type>
<position>-14,-11.5</position>
<output>
<ID>OUT_0</ID>38 </output>
<input>
<ID>clock</ID>36 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>81</ID>
<type>AE_DFF_LOW</type>
<position>11,-12.5</position>
<output>
<ID>OUT_0</ID>39 </output>
<input>
<ID>clock</ID>36 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>82</ID>
<type>AE_DFF_LOW</type>
<position>34.5,-13.5</position>
<output>
<ID>OUT_0</ID>40 </output>
<input>
<ID>clock</ID>36 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_TOGGLE</type>
<position>-58.5,-33</position>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>88</ID>
<type>GA_LED</type>
<position>-38,0</position>
<input>
<ID>N_in2</ID>37 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>GA_LED</type>
<position>-16,0</position>
<input>
<ID>N_in2</ID>38 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>GA_LED</type>
<position>9,-0.5</position>
<input>
<ID>N_in2</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>GA_LED</type>
<position>32.5,-0.5</position>
<input>
<ID>N_in1</ID>41 </input>
<input>
<ID>N_in2</ID>40 </input>
<input>
<ID>N_in3</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>95</ID>
<type>AA_TOGGLE</type>
<position>-54.5,-35</position>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44,-45.5,-44,-37.5</points>
<connection>
<GID>58</GID>
<name>IN_3</name></connection>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20,-45.5,-20,-38</points>
<connection>
<GID>59</GID>
<name>IN_3</name></connection>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-46,3,-38.5</points>
<connection>
<GID>60</GID>
<name>IN_3</name></connection>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-46,25.5,-39</points>
<connection>
<GID>61</GID>
<name>IN_3</name></connection>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-21.5,35.5,-16.5</points>
<connection>
<GID>82</GID>
<name>clock</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-48.5,-21.5,35.5,-21.5</points>
<intersection>-48.5 7</intersection>
<intersection>-35 4</intersection>
<intersection>-13 5</intersection>
<intersection>12 6</intersection>
<intersection>35.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-35,-21.5,-35,-14</points>
<connection>
<GID>79</GID>
<name>clock</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-13,-21.5,-13,-14.5</points>
<connection>
<GID>80</GID>
<name>clock</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>12,-21.5,12,-15.5</points>
<connection>
<GID>81</GID>
<name>clock</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-48.5,-22.5,-48.5,-21.5</points>
<connection>
<GID>77</GID>
<name>CLK</name></connection>
<intersection>-21.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27,-43.5,-27,-6</points>
<intersection>-43.5 6</intersection>
<intersection>-6 7</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-42,-43.5,-27,-43.5</points>
<intersection>-42 10</intersection>
<intersection>-27 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-38,-6,-27,-6</points>
<intersection>-38 9</intersection>
<intersection>-27 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-38,-8,-38,-1</points>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection>
<connection>
<GID>88</GID>
<name>N_in2</name></connection>
<intersection>-6 7</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-42,-43.5,-42,-37.5</points>
<connection>
<GID>58</GID>
<name>IN_2</name></connection>
<intersection>-43.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-43.5,-6,-6.5</points>
<intersection>-43.5 7</intersection>
<intersection>-6.5 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-18,-43.5,-6,-43.5</points>
<intersection>-18 11</intersection>
<intersection>-6 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-16,-6.5,-6,-6.5</points>
<intersection>-16 10</intersection>
<intersection>-6 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-16,-8.5,-16,-1</points>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection>
<connection>
<GID>90</GID>
<name>N_in2</name></connection>
<intersection>-6.5 8</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-18,-43.5,-18,-38</points>
<connection>
<GID>59</GID>
<name>IN_2</name></connection>
<intersection>-43.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-43,18.5,-7</points>
<intersection>-43 4</intersection>
<intersection>-7 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>5,-43,18.5,-43</points>
<intersection>5 7</intersection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>9,-7,18.5,-7</points>
<intersection>9 8</intersection>
<intersection>18.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>5,-43,5,-38.5</points>
<connection>
<GID>60</GID>
<name>IN_2</name></connection>
<intersection>-43 4</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>9,-9.5,9,-1.5</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<connection>
<GID>92</GID>
<name>N_in2</name></connection>
<intersection>-7 5</intersection></vsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-45.5,42,-7.5</points>
<intersection>-45.5 4</intersection>
<intersection>-7.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>27.5,-45.5,42,-45.5</points>
<intersection>27.5 8</intersection>
<intersection>42 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>32.5,-7.5,42,-7.5</points>
<intersection>32.5 7</intersection>
<intersection>42 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>32.5,-10.5,32.5,-1.5</points>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection>
<connection>
<GID>94</GID>
<name>N_in2</name></connection>
<intersection>-7.5 5</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>27.5,-45.5,27.5,-39</points>
<connection>
<GID>61</GID>
<name>IN_2</name></connection>
<intersection>-45.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-0.5,32.5,0.5</points>
<connection>
<GID>94</GID>
<name>N_in3</name></connection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-0.5,33.5,-0.5</points>
<connection>
<GID>94</GID>
<name>N_in1</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-52.5,-36,23.5,-36</points>
<connection>
<GID>61</GID>
<name>SEL_1</name></connection>
<intersection>-52.5 3</intersection>
<intersection>-46 6</intersection>
<intersection>-22 4</intersection>
<intersection>1 8</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-52.5,-36,-52.5,-35</points>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection>
<intersection>-36 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-22,-36,-22,-35</points>
<connection>
<GID>59</GID>
<name>SEL_1</name></connection>
<intersection>-36 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-46,-36,-46,-34.5</points>
<connection>
<GID>58</GID>
<name>SEL_1</name></connection>
<intersection>-36 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>1,-36,1,-35.5</points>
<connection>
<GID>60</GID>
<name>SEL_1</name></connection>
<intersection>-36 1</intersection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-56.5,-33,-22,-33</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>-46 8</intersection>
<intersection>-22 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-22,-34,-22,-33</points>
<connection>
<GID>59</GID>
<name>SEL_0</name></connection>
<intersection>-33.5 9</intersection>
<intersection>-33 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-46,-33.5,-46,-33</points>
<connection>
<GID>58</GID>
<name>SEL_0</name></connection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-22,-33.5,1,-33.5</points>
<intersection>-22 5</intersection>
<intersection>1 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>1,-34.5,1,-33.5</points>
<connection>
<GID>60</GID>
<name>SEL_0</name></connection>
<intersection>-34 11</intersection>
<intersection>-33.5 9</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>1,-34,23.5,-34</points>
<intersection>1 10</intersection>
<intersection>23.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>23.5,-35,23.5,-34</points>
<connection>
<GID>61</GID>
<name>SEL_0</name></connection>
<intersection>-34 11</intersection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31.5,-39,-31.5,-8</points>
<intersection>-39 3</intersection>
<intersection>-8 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-38,-39,-16,-39</points>
<intersection>-38 5</intersection>
<intersection>-31.5 0</intersection>
<intersection>-16 11</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-35,-8,-31.5,-8</points>
<connection>
<GID>79</GID>
<name>OUTINV_0</name></connection>
<intersection>-31.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-38,-39,-38,-37.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>-39 3</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-16,-39,-16,-38</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>-39 3</intersection></vsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-39.5,29.5,-39</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>-39.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>9,-39.5,29.5,-39.5</points>
<intersection>9 3</intersection>
<intersection>29.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>9,-39.5,9,-38.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>-39.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-39.5,7,-38.5</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>-39.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-14,-39.5,7,-39.5</points>
<intersection>-14 3</intersection>
<intersection>7 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-14,-39.5,-14,-38</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>-39.5 2</intersection></vsegment></shape></wire></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>