<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>36.5,-39.9583,84.5,-63.6838</PageViewport>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>52.5,-25.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>43.5,-24</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>43.5,-27</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>59,-25.5</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>50,-20.5</position>
<gparam>LABEL_TEXT AND Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>39.5,-24</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>39.5,-27</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>63.5,-25</position>
<gparam>LABEL_TEXT Y = A.B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>75.5,-20.5</position>
<gparam>LABEL_TEXT Truth Table</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>74.5,-23.5</position>
<gparam>LABEL_TEXT A    B    Y</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>74.5,-25</position>
<gparam>LABEL_TEXT 0    0    0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>74.5,-26.5</position>
<gparam>LABEL_TEXT 0    1    0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>74.5,-28</position>
<gparam>LABEL_TEXT 1    0    0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>74.5,-29.5</position>
<gparam>LABEL_TEXT 1    1    1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>49,-32.5</position>
<gparam>LABEL_TEXT OR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_TOGGLE</type>
<position>43.5,-37</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>43.5,-40</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>33</ID>
<type>GA_LED</type>
<position>59,-38.5</position>
<input>
<ID>N_in0</ID>6 </input>
<input>
<ID>N_in2</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>39.5,-37</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>39.5,-40</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>63.5,-38</position>
<gparam>LABEL_TEXT Y = A+B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AE_OR2</type>
<position>52.5,-38.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>50,-45.5</position>
<gparam>LABEL_TEXT NOT Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_INVERTER</type>
<position>54,-50</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_TOGGLE</type>
<position>44,-50</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>44</ID>
<type>GA_LED</type>
<position>61,-50</position>
<input>
<ID>N_in0</ID>8 </input>
<input>
<ID>N_in1</ID>8 </input>
<input>
<ID>N_in3</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>64.5,-50</position>
<gparam>LABEL_TEXT Y = A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>66,-48.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>51,-55.5</position>
<gparam>LABEL_TEXT NAND Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>AA_LABEL</type>
<position>50,-68</position>
<gparam>LABEL_TEXT NOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>51.5,-79</position>
<gparam>LABEL_TEXT X-NOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>51.5,-91</position>
<gparam>LABEL_TEXT X-OR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AO_XNOR2</type>
<position>52.5,-86.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>58</ID>
<type>AI_XOR2</type>
<position>54.5,-97</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>60</ID>
<type>BA_NAND2</type>
<position>51,-62</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>62</ID>
<type>BE_NOR2</type>
<position>52,-74</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_TOGGLE</type>
<position>41.5,-60.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>65</ID>
<type>AA_TOGGLE</type>
<position>41.5,-63.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>61.5,-61.5</position>
<gparam>LABEL_TEXT Y = A.B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_TOGGLE</type>
<position>42,-73</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_TOGGLE</type>
<position>42,-76</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>62,-74</position>
<gparam>LABEL_TEXT Y = A+B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_TOGGLE</type>
<position>39.5,-96</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>71</ID>
<type>AA_TOGGLE</type>
<position>39.5,-99</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_TOGGLE</type>
<position>41,-85</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_TOGGLE</type>
<position>41,-88</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_LABEL</type>
<position>65.5,-86.5</position>
<gparam>LABEL_TEXT Y = A.B + A.B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>GA_LED</type>
<position>57.5,-62</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>GA_LED</type>
<position>57,-74</position>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>GA_LED</type>
<position>59.5,-97</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>GA_LED</type>
<position>58,-86.5</position>
<input>
<ID>N_in0</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>63,-60</position>
<gparam>LABEL_TEXT ___</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>63.5,-72.5</position>
<gparam>LABEL_TEXT ____</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>64,-85</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>70,-85</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_LABEL</type>
<position>66.5,-97</position>
<gparam>LABEL_TEXT Y = A.B + A.B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>AA_LABEL</type>
<position>65,-95.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>AA_LABEL</type>
<position>66.5,-95.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-24,49.5,-24</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>49.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>49.5,-24.5,49.5,-24</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-24 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-27,49.5,-27</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>49.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>49.5,-27,49.5,-26.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-27 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55.5,-25.5,58,-25.5</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>8</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-37.5,47.5,-37</points>
<intersection>-37.5 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-37.5,49.5,-37.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-37,47.5,-37</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-40,47.5,-39.5</points>
<intersection>-40 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-39.5,49.5,-39.5</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-40,47.5,-40</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55.5,-38.5,59,-38.5</points>
<connection>
<GID>33</GID>
<name>N_in0</name></connection>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>59 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>59,-39.5,59,-38.5</points>
<connection>
<GID>33</GID>
<name>N_in2</name></connection>
<intersection>-38.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46,-50,51,-50</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<connection>
<GID>42</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-50,62,-50</points>
<connection>
<GID>44</GID>
<name>N_in1</name></connection>
<connection>
<GID>44</GID>
<name>N_in0</name></connection>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>61 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>61,-50,61,-49</points>
<connection>
<GID>44</GID>
<name>N_in3</name></connection>
<intersection>-50 1</intersection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-61,45.5,-60.5</points>
<intersection>-61 1</intersection>
<intersection>-60.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,-61,48,-61</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>45.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-60.5,45.5,-60.5</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-63.5,45.5,-63</points>
<intersection>-63.5 2</intersection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,-63,48,-63</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>45.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-63.5,45.5,-63.5</points>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-62,56.5,-62</points>
<connection>
<GID>80</GID>
<name>N_in0</name></connection>
<connection>
<GID>60</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-73,49,-73</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-76,46.5,-75</points>
<intersection>-76 2</intersection>
<intersection>-75 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-75,49,-75</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>44,-76,46.5,-76</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41.5,-96,51.5,-96</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-98.5,46.5,-98</points>
<intersection>-98.5 2</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-98,51.5,-98</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-98.5,51,-98.5</points>
<intersection>46.5 0</intersection>
<intersection>51 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>51,-99,51,-98.5</points>
<intersection>-99 4</intersection>
<intersection>-98.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>41.5,-99,51,-99</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<intersection>51 3</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57.5,-97,58.5,-97</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<connection>
<GID>84</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-85.5,46.5,-85</points>
<intersection>-85.5 1</intersection>
<intersection>-85 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-85.5,49.5,-85.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43,-85,46.5,-85</points>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-88,46.5,-87.5</points>
<intersection>-88 2</intersection>
<intersection>-87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-87.5,49.5,-87.5</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43,-88,46.5,-88</points>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55.5,-86.5,57,-86.5</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<connection>
<GID>86</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-216.283,57.3852,73.85,-86.0222</PageViewport>
<gate>
<ID>193</ID>
<type>AA_LABEL</type>
<position>112,31.5</position>
<gparam>LABEL_TEXT NAND Gate as UNIVERSAL GATE</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>194</ID>
<type>BA_NAND2</type>
<position>57.5,0</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>195</ID>
<type>BA_NAND2</type>
<position>72,0</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>78 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>196</ID>
<type>GA_LED</type>
<position>79,0</position>
<input>
<ID>N_in0</ID>79 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>197</ID>
<type>AA_LABEL</type>
<position>86,0.5</position>
<gparam>LABEL_TEXT Output Y=A.B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>198</ID>
<type>AA_TOGGLE</type>
<position>47.5,1</position>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>199</ID>
<type>AA_LABEL</type>
<position>41,1.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>200</ID>
<type>AA_TOGGLE</type>
<position>47.5,-2</position>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>201</ID>
<type>AA_LABEL</type>
<position>41.5,-2</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>202</ID>
<type>AA_LABEL</type>
<position>63.5,6.5</position>
<gparam>LABEL_TEXT NAND as AND Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>203</ID>
<type>BA_NAND2</type>
<position>56.5,-19.5</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>204</ID>
<type>BA_NAND2</type>
<position>56.5,-26.5</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>83 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>205</ID>
<type>GA_LED</type>
<position>78,-19.5</position>
<input>
<ID>N_in0</ID>86 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>206</ID>
<type>AA_LABEL</type>
<position>85,-19</position>
<gparam>LABEL_TEXT Output Y=A.B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>207</ID>
<type>AA_TOGGLE</type>
<position>46.5,-18.5</position>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>208</ID>
<type>AA_LABEL</type>
<position>40,-18</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>209</ID>
<type>AA_TOGGLE</type>
<position>46.5,-27</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>210</ID>
<type>AA_LABEL</type>
<position>41,-27</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>211</ID>
<type>AA_LABEL</type>
<position>63.5,-11.5</position>
<gparam>LABEL_TEXT NAND as OR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>212</ID>
<type>BA_NAND2</type>
<position>67.5,-22</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>213</ID>
<type>BA_NAND2</type>
<position>54.5,-44</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>214</ID>
<type>BA_NAND2</type>
<position>54.5,-51</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>88 </input>
<output>
<ID>OUT</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>215</ID>
<type>GA_LED</type>
<position>77.5,-46.5</position>
<input>
<ID>N_in0</ID>91 </input>
<input>
<ID>N_in1</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>216</ID>
<type>AA_LABEL</type>
<position>91,-46</position>
<gparam>LABEL_TEXT Output Y=(A+B)'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>217</ID>
<type>AA_TOGGLE</type>
<position>44.5,-43</position>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>218</ID>
<type>AA_LABEL</type>
<position>38,-42.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>219</ID>
<type>AA_TOGGLE</type>
<position>44.5,-51.5</position>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>220</ID>
<type>AA_LABEL</type>
<position>39,-51.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>221</ID>
<type>AA_LABEL</type>
<position>61.5,-36</position>
<gparam>LABEL_TEXT NAND as NOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>222</ID>
<type>BA_NAND2</type>
<position>65.5,-46.5</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>223</ID>
<type>BA_NAND2</type>
<position>72.5,-46.5</position>
<input>
<ID>IN_0</ID>92 </input>
<input>
<ID>IN_1</ID>92 </input>
<output>
<ID>OUT</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>224</ID>
<type>GA_LED</type>
<position>164.5,14.5</position>
<input>
<ID>N_in0</ID>98 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>225</ID>
<type>AA_LABEL</type>
<position>173.5,15</position>
<gparam>LABEL_TEXT Output Y=A'B+AB'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>226</ID>
<type>AA_TOGGLE</type>
<position>133,15.5</position>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>227</ID>
<type>AA_LABEL</type>
<position>126.5,16</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>228</ID>
<type>AA_TOGGLE</type>
<position>133,7</position>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>229</ID>
<type>AA_LABEL</type>
<position>127.5,7</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>230</ID>
<type>AA_LABEL</type>
<position>150,22.5</position>
<gparam>LABEL_TEXT NAND as XOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>231</ID>
<type>BA_NAND2</type>
<position>143,11.5</position>
<input>
<ID>IN_0</ID>93 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>232</ID>
<type>BA_NAND2</type>
<position>153,15.5</position>
<input>
<ID>IN_0</ID>93 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>233</ID>
<type>BA_NAND2</type>
<position>152.5,7.5</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>234</ID>
<type>BA_NAND2</type>
<position>159.5,12</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>235</ID>
<type>GA_LED</type>
<position>176,-25</position>
<input>
<ID>N_in0</ID>105 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>236</ID>
<type>AA_LABEL</type>
<position>185,-24.5</position>
<gparam>LABEL_TEXT Output Y=A'B+AB'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>237</ID>
<type>AA_TOGGLE</type>
<position>133.5,-21.5</position>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>238</ID>
<type>AA_LABEL</type>
<position>127,-21</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>239</ID>
<type>AA_TOGGLE</type>
<position>133.5,-30</position>
<output>
<ID>OUT_0</ID>100 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>240</ID>
<type>AA_LABEL</type>
<position>128,-30</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>241</ID>
<type>AA_LABEL</type>
<position>150.5,-14.5</position>
<gparam>LABEL_TEXT NAND as XNOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>242</ID>
<type>BA_NAND2</type>
<position>143.5,-25.5</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>100 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>243</ID>
<type>BA_NAND2</type>
<position>153.5,-21.5</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>101 </input>
<output>
<ID>OUT</ID>102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>244</ID>
<type>BA_NAND2</type>
<position>153,-29.5</position>
<input>
<ID>IN_0</ID>101 </input>
<input>
<ID>IN_1</ID>100 </input>
<output>
<ID>OUT</ID>103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>245</ID>
<type>BA_NAND2</type>
<position>160,-25</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>103 </input>
<output>
<ID>OUT</ID>104 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>246</ID>
<type>BA_NAND2</type>
<position>168,-25</position>
<input>
<ID>IN_0</ID>104 </input>
<input>
<ID>IN_1</ID>104 </input>
<output>
<ID>OUT</ID>105 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>247</ID>
<type>GA_LED</type>
<position>-119.5,-48.5</position>
<input>
<ID>N_in0</ID>122 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>248</ID>
<type>AA_TOGGLE</type>
<position>-161.5,12</position>
<output>
<ID>OUT_0</ID>109 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>249</ID>
<type>GA_LED</type>
<position>-139,12.5</position>
<input>
<ID>N_in0</ID>108 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>250</ID>
<type>AA_LABEL</type>
<position>-168,12.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>251</ID>
<type>AA_LABEL</type>
<position>-132,13</position>
<gparam>LABEL_TEXT Output Y=A'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>252</ID>
<type>AA_LABEL</type>
<position>-147.5,19.5</position>
<gparam>LABEL_TEXT NOR as NOT Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>253</ID>
<type>AA_LABEL</type>
<position>-112.5,-48</position>
<gparam>LABEL_TEXT Output Y=(A.B)'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>254</ID>
<type>GA_LED</type>
<position>-132,-3.5</position>
<input>
<ID>N_in0</ID>112 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>255</ID>
<type>AA_LABEL</type>
<position>-125,-3</position>
<gparam>LABEL_TEXT Output Y=A+B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>256</ID>
<type>AA_TOGGLE</type>
<position>-163.5,-2.5</position>
<output>
<ID>OUT_0</ID>114 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>257</ID>
<type>AA_LABEL</type>
<position>-170,-2</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>258</ID>
<type>AA_TOGGLE</type>
<position>-163.5,-5.5</position>
<output>
<ID>OUT_0</ID>113 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>259</ID>
<type>BE_NOR2</type>
<position>-150,12.5</position>
<input>
<ID>IN_0</ID>109 </input>
<input>
<ID>IN_1</ID>109 </input>
<output>
<ID>OUT</ID>108 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>260</ID>
<type>AA_LABEL</type>
<position>-169.5,-5.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>261</ID>
<type>AA_LABEL</type>
<position>-147.5,3</position>
<gparam>LABEL_TEXT NOR as OR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>262</ID>
<type>GA_LED</type>
<position>-128,-24</position>
<input>
<ID>N_in0</ID>118 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>263</ID>
<type>BE_NOR2</type>
<position>-154,-4</position>
<input>
<ID>IN_0</ID>114 </input>
<input>
<ID>IN_1</ID>113 </input>
<output>
<ID>OUT</ID>111 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>264</ID>
<type>AA_LABEL</type>
<position>-121,-23.5</position>
<gparam>LABEL_TEXT Output Y=A.B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>265</ID>
<type>BE_NOR2</type>
<position>-140.5,-4</position>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>111 </input>
<output>
<ID>OUT</ID>112 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>266</ID>
<type>AA_TOGGLE</type>
<position>-160.5,-20.5</position>
<output>
<ID>OUT_0</ID>120 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>267</ID>
<type>AA_LABEL</type>
<position>-167,-20</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>268</ID>
<type>AA_TOGGLE</type>
<position>-160.5,-29</position>
<output>
<ID>OUT_0</ID>119 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>269</ID>
<type>AA_LABEL</type>
<position>-166,-29</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>270</ID>
<type>AA_LABEL</type>
<position>-143.5,-13.5</position>
<gparam>LABEL_TEXT NOR as AND Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>271</ID>
<type>AA_TOGGLE</type>
<position>-159.5,-44</position>
<output>
<ID>OUT_0</ID>115 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>272</ID>
<type>AA_LABEL</type>
<position>-166,-43.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>273</ID>
<type>BE_NOR2</type>
<position>-151,-20.5</position>
<input>
<ID>IN_0</ID>120 </input>
<input>
<ID>IN_1</ID>120 </input>
<output>
<ID>OUT</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>274</ID>
<type>AA_TOGGLE</type>
<position>-159.5,-52.5</position>
<output>
<ID>OUT_0</ID>110 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>275</ID>
<type>BE_NOR2</type>
<position>-151,-29</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>117 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>276</ID>
<type>AA_LABEL</type>
<position>-165,-52.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>277</ID>
<type>BE_NOR2</type>
<position>-138,-25</position>
<input>
<ID>IN_0</ID>116 </input>
<input>
<ID>IN_1</ID>117 </input>
<output>
<ID>OUT</ID>118 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>278</ID>
<type>AA_LABEL</type>
<position>-142.5,-37</position>
<gparam>LABEL_TEXT NOR as NAND Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>279</ID>
<type>BE_NOR2</type>
<position>-150,-44</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>115 </input>
<output>
<ID>OUT</ID>106 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>280</ID>
<type>BE_NOR2</type>
<position>-150,-52.5</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>110 </input>
<output>
<ID>OUT</ID>107 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>281</ID>
<type>BE_NOR2</type>
<position>-137,-48.5</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>107 </input>
<output>
<ID>OUT</ID>121 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>282</ID>
<type>GA_LED</type>
<position>-40.5,14</position>
<input>
<ID>N_in0</ID>123 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>283</ID>
<type>BE_NOR2</type>
<position>-128,-48.5</position>
<input>
<ID>IN_0</ID>121 </input>
<input>
<ID>IN_1</ID>121 </input>
<output>
<ID>OUT</ID>122 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>284</ID>
<type>AA_LABEL</type>
<position>-31.5,14.5</position>
<gparam>LABEL_TEXT Output Y=A'B+AB'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>285</ID>
<type>AA_TOGGLE</type>
<position>-83,17.5</position>
<output>
<ID>OUT_0</ID>125 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>286</ID>
<type>AA_LABEL</type>
<position>-89.5,18</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>287</ID>
<type>AA_TOGGLE</type>
<position>-83,9</position>
<output>
<ID>OUT_0</ID>124 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>288</ID>
<type>AA_LABEL</type>
<position>-88.5,9</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>289</ID>
<type>AA_LABEL</type>
<position>-66,24.5</position>
<gparam>LABEL_TEXT NAND as XOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>290</ID>
<type>BE_NOR2</type>
<position>-71.5,13.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>124 </input>
<output>
<ID>OUT</ID>126 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>291</ID>
<type>BE_NOR2</type>
<position>-60.5,17</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>126 </input>
<output>
<ID>OUT</ID>127 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>292</ID>
<type>BE_NOR2</type>
<position>-60.5,8.5</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>124 </input>
<output>
<ID>OUT</ID>128 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>293</ID>
<type>BE_NOR2</type>
<position>-53.5,13</position>
<input>
<ID>IN_0</ID>127 </input>
<input>
<ID>IN_1</ID>128 </input>
<output>
<ID>OUT</ID>129 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>294</ID>
<type>BE_NOR2</type>
<position>-46.5,13</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>129 </input>
<output>
<ID>OUT</ID>123 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>295</ID>
<type>GA_LED</type>
<position>-26,-17.5</position>
<input>
<ID>N_in0</ID>137 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>296</ID>
<type>AA_LABEL</type>
<position>-17,-17</position>
<gparam>LABEL_TEXT Output Y=AB+A'B'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>297</ID>
<type>AA_TOGGLE</type>
<position>-85.5,-13</position>
<output>
<ID>OUT_0</ID>131 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>298</ID>
<type>AA_LABEL</type>
<position>-92,-12.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>299</ID>
<type>AA_TOGGLE</type>
<position>-85.5,-21.5</position>
<output>
<ID>OUT_0</ID>130 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>300</ID>
<type>AA_LABEL</type>
<position>-91,-21.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>301</ID>
<type>AA_LABEL</type>
<position>-68.5,-6</position>
<gparam>LABEL_TEXT NAND as XNOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>302</ID>
<type>BE_NOR2</type>
<position>-74,-17</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>132 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>303</ID>
<type>BE_NOR2</type>
<position>-63,-13.5</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>132 </input>
<output>
<ID>OUT</ID>133 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>304</ID>
<type>BE_NOR2</type>
<position>-63,-22</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>305</ID>
<type>BE_NOR2</type>
<position>-56,-17.5</position>
<input>
<ID>IN_0</ID>133 </input>
<input>
<ID>IN_1</ID>134 </input>
<output>
<ID>OUT</ID>135 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>306</ID>
<type>BE_NOR2</type>
<position>-49,-17.5</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>135 </input>
<output>
<ID>OUT</ID>136 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>307</ID>
<type>BE_NOR2</type>
<position>-39.5,-17.5</position>
<input>
<ID>IN_0</ID>136 </input>
<input>
<ID>IN_1</ID>136 </input>
<output>
<ID>OUT</ID>137 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>308</ID>
<type>AA_LABEL</type>
<position>-111,34.5</position>
<gparam>LABEL_TEXT NOR as UNIVERSAL GATES</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>187</ID>
<type>BA_NAND2</type>
<position>63.5,14</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_1</ID>76 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>188</ID>
<type>AA_TOGGLE</type>
<position>49,13.5</position>
<output>
<ID>OUT_0</ID>76 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>189</ID>
<type>GA_LED</type>
<position>71.5,14</position>
<input>
<ID>N_in0</ID>77 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>190</ID>
<type>AA_LABEL</type>
<position>42.5,14</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>191</ID>
<type>AA_LABEL</type>
<position>78.5,14.5</position>
<gparam>LABEL_TEXT Output Y=A'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>192</ID>
<type>AA_LABEL</type>
<position>63,21</position>
<gparam>LABEL_TEXT NAND as NOT Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51,13.5,60.5,13.5</points>
<connection>
<GID>188</GID>
<name>OUT_0</name></connection>
<intersection>60.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>60.5,13,60.5,15</points>
<connection>
<GID>187</GID>
<name>IN_1</name></connection>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>13.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>66.5,14,70.5,14</points>
<connection>
<GID>187</GID>
<name>OUT</name></connection>
<connection>
<GID>189</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-1,69,1</points>
<connection>
<GID>195</GID>
<name>IN_1</name></connection>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,0,69,0</points>
<connection>
<GID>194</GID>
<name>OUT</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,0,78,0</points>
<connection>
<GID>195</GID>
<name>OUT</name></connection>
<connection>
<GID>196</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,1,54.5,1</points>
<connection>
<GID>198</GID>
<name>OUT_0</name></connection>
<connection>
<GID>194</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-2,52,-1</points>
<intersection>-2 2</intersection>
<intersection>-1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-1,54.5,-1</points>
<connection>
<GID>194</GID>
<name>IN_1</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-2,52,-2</points>
<connection>
<GID>200</GID>
<name>OUT_0</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-20.5,53.5,-18.5</points>
<connection>
<GID>203</GID>
<name>IN_1</name></connection>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48.5,-18.5,53.5,-18.5</points>
<connection>
<GID>207</GID>
<name>OUT_0</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-27.5,53.5,-25.5</points>
<connection>
<GID>204</GID>
<name>IN_1</name></connection>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48.5,-27,53.5,-27</points>
<connection>
<GID>209</GID>
<name>OUT_0</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-26.5,62,-23</points>
<intersection>-26.5 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-23,64.5,-23</points>
<connection>
<GID>212</GID>
<name>IN_1</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59.5,-26.5,62,-26.5</points>
<connection>
<GID>204</GID>
<name>OUT</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-21,62,-19.5</points>
<intersection>-21 1</intersection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-21,64.5,-21</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59.5,-19.5,62,-19.5</points>
<connection>
<GID>203</GID>
<name>OUT</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-22,73.5,-19.5</points>
<intersection>-22 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-19.5,77,-19.5</points>
<connection>
<GID>205</GID>
<name>N_in0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-22,73.5,-22</points>
<connection>
<GID>212</GID>
<name>OUT</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-45,51.5,-43</points>
<connection>
<GID>213</GID>
<name>IN_1</name></connection>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-43,51.5,-43</points>
<connection>
<GID>217</GID>
<name>OUT_0</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-52,51.5,-50</points>
<connection>
<GID>214</GID>
<name>IN_1</name></connection>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-51.5,51.5,-51.5</points>
<connection>
<GID>219</GID>
<name>OUT_0</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-51,60,-47.5</points>
<intersection>-51 2</intersection>
<intersection>-47.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60,-47.5,62.5,-47.5</points>
<connection>
<GID>222</GID>
<name>IN_1</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-51,60,-51</points>
<connection>
<GID>214</GID>
<name>OUT</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-45.5,60,-44</points>
<intersection>-45.5 1</intersection>
<intersection>-44 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60,-45.5,62.5,-45.5</points>
<connection>
<GID>222</GID>
<name>IN_0</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-44,60,-44</points>
<connection>
<GID>213</GID>
<name>OUT</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75.5,-46.5,78.5,-46.5</points>
<connection>
<GID>223</GID>
<name>OUT</name></connection>
<connection>
<GID>215</GID>
<name>N_in0</name></connection>
<connection>
<GID>215</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-47.5,69.5,-45.5</points>
<connection>
<GID>223</GID>
<name>IN_1</name></connection>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-46.5,69.5,-46.5</points>
<connection>
<GID>222</GID>
<name>OUT</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,15.5,142.5,16.5</points>
<intersection>15.5 2</intersection>
<intersection>16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142.5,16.5,150,16.5</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>135,15.5,142.5,15.5</points>
<connection>
<GID>226</GID>
<name>OUT_0</name></connection>
<intersection>140 3</intersection>
<intersection>142.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>140,12.5,140,15.5</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>15.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,6.5,142,7</points>
<intersection>6.5 1</intersection>
<intersection>7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142,6.5,149.5,6.5</points>
<connection>
<GID>233</GID>
<name>IN_1</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>135,7,142,7</points>
<connection>
<GID>228</GID>
<name>OUT_0</name></connection>
<intersection>140 3</intersection>
<intersection>142 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>140,7,140,10.5</points>
<connection>
<GID>231</GID>
<name>IN_1</name></connection>
<intersection>7 2</intersection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147.5,8.5,147.5,14.5</points>
<intersection>8.5 1</intersection>
<intersection>11.5 2</intersection>
<intersection>14.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147.5,8.5,149.5,8.5</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>147.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>146,11.5,147.5,11.5</points>
<connection>
<GID>231</GID>
<name>OUT</name></connection>
<intersection>147.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>147.5,14.5,150,14.5</points>
<connection>
<GID>232</GID>
<name>IN_1</name></connection>
<intersection>147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,13,156,15.5</points>
<connection>
<GID>232</GID>
<name>OUT</name></connection>
<intersection>13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156,13,156.5,13</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,7.5,156,11</points>
<intersection>7.5 2</intersection>
<intersection>11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156,11,156.5,11</points>
<connection>
<GID>234</GID>
<name>IN_1</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155.5,7.5,156,7.5</points>
<connection>
<GID>233</GID>
<name>OUT</name></connection>
<intersection>156 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,12,163,14.5</points>
<intersection>12 2</intersection>
<intersection>14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>163,14.5,163.5,14.5</points>
<connection>
<GID>224</GID>
<name>N_in0</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162.5,12,163,12</points>
<connection>
<GID>234</GID>
<name>OUT</name></connection>
<intersection>163 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,-21.5,143,-20.5</points>
<intersection>-21.5 2</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143,-20.5,150.5,-20.5</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>143 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>135.5,-21.5,143,-21.5</points>
<connection>
<GID>237</GID>
<name>OUT_0</name></connection>
<intersection>140.5 3</intersection>
<intersection>143 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>140.5,-24.5,140.5,-21.5</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>-21.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-30.5,142.5,-30</points>
<intersection>-30.5 1</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142.5,-30.5,150,-30.5</points>
<connection>
<GID>244</GID>
<name>IN_1</name></connection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>135.5,-30,142.5,-30</points>
<connection>
<GID>239</GID>
<name>OUT_0</name></connection>
<intersection>140.5 3</intersection>
<intersection>142.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>140.5,-30,140.5,-26.5</points>
<connection>
<GID>242</GID>
<name>IN_1</name></connection>
<intersection>-30 2</intersection></vsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148,-28.5,148,-22.5</points>
<intersection>-28.5 1</intersection>
<intersection>-25.5 2</intersection>
<intersection>-22.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>148,-28.5,150,-28.5</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>148 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>146.5,-25.5,148,-25.5</points>
<connection>
<GID>242</GID>
<name>OUT</name></connection>
<intersection>148 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>148,-22.5,150.5,-22.5</points>
<connection>
<GID>243</GID>
<name>IN_1</name></connection>
<intersection>148 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-24,156.5,-21.5</points>
<connection>
<GID>243</GID>
<name>OUT</name></connection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156.5,-24,157,-24</points>
<connection>
<GID>245</GID>
<name>IN_0</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-29.5,156.5,-26</points>
<intersection>-29.5 2</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156.5,-26,157,-26</points>
<connection>
<GID>245</GID>
<name>IN_1</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156,-29.5,156.5,-29.5</points>
<connection>
<GID>244</GID>
<name>OUT</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>163,-25,165,-25</points>
<connection>
<GID>245</GID>
<name>OUT</name></connection>
<intersection>165 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>165,-26,165,-24</points>
<connection>
<GID>246</GID>
<name>IN_1</name></connection>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<intersection>-25 1</intersection></vsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>171,-25,175,-25</points>
<connection>
<GID>246</GID>
<name>OUT</name></connection>
<connection>
<GID>235</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-143.5,-47.5,-143.5,-44</points>
<intersection>-47.5 1</intersection>
<intersection>-44 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-143.5,-47.5,-140,-47.5</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>-143.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-147,-44,-143.5,-44</points>
<connection>
<GID>279</GID>
<name>OUT</name></connection>
<intersection>-143.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-143.5,-52.5,-143.5,-49.5</points>
<intersection>-52.5 2</intersection>
<intersection>-49.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-143.5,-49.5,-140,-49.5</points>
<connection>
<GID>281</GID>
<name>IN_1</name></connection>
<intersection>-143.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-147,-52.5,-143.5,-52.5</points>
<connection>
<GID>280</GID>
<name>OUT</name></connection>
<intersection>-143.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-147,12.5,-140,12.5</points>
<connection>
<GID>259</GID>
<name>OUT</name></connection>
<connection>
<GID>249</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-153,11.5,-153,13.5</points>
<connection>
<GID>259</GID>
<name>IN_1</name></connection>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<intersection>12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-159.5,12,-153,12</points>
<connection>
<GID>248</GID>
<name>OUT_0</name></connection>
<intersection>-153 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-153,-53.5,-153,-51.5</points>
<connection>
<GID>280</GID>
<name>IN_1</name></connection>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-157.5,-52.5,-153,-52.5</points>
<connection>
<GID>274</GID>
<name>OUT_0</name></connection>
<intersection>-153 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-143.5,-5,-143.5,-3</points>
<connection>
<GID>265</GID>
<name>IN_1</name></connection>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<intersection>-4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-151,-4,-143.5,-4</points>
<connection>
<GID>263</GID>
<name>OUT</name></connection>
<intersection>-143.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-135.5,-4,-135.5,-3.5</points>
<intersection>-4 2</intersection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-135.5,-3.5,-133,-3.5</points>
<connection>
<GID>254</GID>
<name>N_in0</name></connection>
<intersection>-135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-137.5,-4,-135.5,-4</points>
<connection>
<GID>265</GID>
<name>OUT</name></connection>
<intersection>-135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-159.5,-5.5,-159.5,-5</points>
<intersection>-5.5 2</intersection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-159.5,-5,-157,-5</points>
<connection>
<GID>263</GID>
<name>IN_1</name></connection>
<intersection>-159.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-161.5,-5.5,-159.5,-5.5</points>
<connection>
<GID>258</GID>
<name>OUT_0</name></connection>
<intersection>-159.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-159.5,-3,-159.5,-2.5</points>
<intersection>-3 1</intersection>
<intersection>-2.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-159.5,-3,-157,-3</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<intersection>-159.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-161.5,-2.5,-159.5,-2.5</points>
<connection>
<GID>256</GID>
<name>OUT_0</name></connection>
<intersection>-159.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-153,-45,-153,-43</points>
<connection>
<GID>279</GID>
<name>IN_1</name></connection>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-157.5,-44,-153,-44</points>
<connection>
<GID>271</GID>
<name>OUT_0</name></connection>
<intersection>-153 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-144.5,-24,-144.5,-20.5</points>
<intersection>-24 1</intersection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-144.5,-24,-141,-24</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>-144.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-148,-20.5,-144.5,-20.5</points>
<connection>
<GID>273</GID>
<name>OUT</name></connection>
<intersection>-144.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-144.5,-29,-144.5,-26</points>
<intersection>-29 2</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-144.5,-26,-141,-26</points>
<connection>
<GID>277</GID>
<name>IN_1</name></connection>
<intersection>-144.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-148,-29,-144.5,-29</points>
<connection>
<GID>275</GID>
<name>OUT</name></connection>
<intersection>-144.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-132,-25,-132,-24</points>
<intersection>-25 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-132,-24,-129,-24</points>
<connection>
<GID>262</GID>
<name>N_in0</name></connection>
<intersection>-132 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-135,-25,-132,-25</points>
<connection>
<GID>277</GID>
<name>OUT</name></connection>
<intersection>-132 0</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-154,-30,-154,-28</points>
<connection>
<GID>275</GID>
<name>IN_1</name></connection>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-158.5,-29,-154,-29</points>
<connection>
<GID>268</GID>
<name>OUT_0</name></connection>
<intersection>-154 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-154,-21.5,-154,-19.5</points>
<connection>
<GID>273</GID>
<name>IN_1</name></connection>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-158.5,-20.5,-154,-20.5</points>
<connection>
<GID>266</GID>
<name>OUT_0</name></connection>
<intersection>-154 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-132.5,-49.5,-132.5,-47.5</points>
<intersection>-49.5 2</intersection>
<intersection>-48.5 1</intersection>
<intersection>-47.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-134,-48.5,-132.5,-48.5</points>
<connection>
<GID>281</GID>
<name>OUT</name></connection>
<intersection>-132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-132.5,-49.5,-131,-49.5</points>
<connection>
<GID>283</GID>
<name>IN_1</name></connection>
<intersection>-132.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-132.5,-47.5,-131,-47.5</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<intersection>-132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-125,-48.5,-120.5,-48.5</points>
<connection>
<GID>283</GID>
<name>OUT</name></connection>
<connection>
<GID>247</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,13,-42.5,14</points>
<intersection>13 2</intersection>
<intersection>14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-42.5,14,-41.5,14</points>
<connection>
<GID>282</GID>
<name>N_in0</name></connection>
<intersection>-42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-43.5,13,-42.5,13</points>
<connection>
<GID>294</GID>
<name>OUT</name></connection>
<intersection>-42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78,7.5,-78,9</points>
<intersection>7.5 1</intersection>
<intersection>9 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-78,7.5,-63.5,7.5</points>
<connection>
<GID>292</GID>
<name>IN_1</name></connection>
<intersection>-78 0</intersection>
<intersection>-74.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-81,9,-78,9</points>
<connection>
<GID>287</GID>
<name>OUT_0</name></connection>
<intersection>-78 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-74.5,7.5,-74.5,12.5</points>
<connection>
<GID>290</GID>
<name>IN_1</name></connection>
<intersection>7.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-81,17.5,-63.5,17.5</points>
<connection>
<GID>285</GID>
<name>OUT_0</name></connection>
<intersection>-74.5 4</intersection>
<intersection>-63.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-63.5,17.5,-63.5,18</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<intersection>17.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-74.5,14.5,-74.5,17.5</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>17.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66,9.5,-66,16</points>
<intersection>9.5 3</intersection>
<intersection>13.5 1</intersection>
<intersection>16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68.5,13.5,-66,13.5</points>
<connection>
<GID>290</GID>
<name>OUT</name></connection>
<intersection>-66 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-66,16,-63.5,16</points>
<connection>
<GID>291</GID>
<name>IN_1</name></connection>
<intersection>-66 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-66,9.5,-63.5,9.5</points>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<intersection>-66 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57,14,-57,17</points>
<intersection>14 1</intersection>
<intersection>17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-57,14,-56.5,14</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>-57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57.5,17,-57,17</points>
<connection>
<GID>291</GID>
<name>OUT</name></connection>
<intersection>-57 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57,8.5,-57,12</points>
<intersection>8.5 2</intersection>
<intersection>12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-57,12,-56.5,12</points>
<connection>
<GID>293</GID>
<name>IN_1</name></connection>
<intersection>-57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57.5,8.5,-57,8.5</points>
<connection>
<GID>292</GID>
<name>OUT</name></connection>
<intersection>-57 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-50,12,-50,14</points>
<intersection>12 3</intersection>
<intersection>13 2</intersection>
<intersection>14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-50,14,-49.5,14</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>-50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-50.5,13,-50,13</points>
<connection>
<GID>293</GID>
<name>OUT</name></connection>
<intersection>-50 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-50,12,-49.5,12</points>
<connection>
<GID>294</GID>
<name>IN_1</name></connection>
<intersection>-50 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-80.5,-23,-80.5,-21.5</points>
<intersection>-23 1</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-80.5,-23,-66,-23</points>
<connection>
<GID>304</GID>
<name>IN_1</name></connection>
<intersection>-80.5 0</intersection>
<intersection>-77 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-83.5,-21.5,-80.5,-21.5</points>
<connection>
<GID>299</GID>
<name>OUT_0</name></connection>
<intersection>-80.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-77,-23,-77,-18</points>
<connection>
<GID>302</GID>
<name>IN_1</name></connection>
<intersection>-23 1</intersection></vsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-83.5,-13,-66,-13</points>
<connection>
<GID>297</GID>
<name>OUT_0</name></connection>
<intersection>-77 4</intersection>
<intersection>-66 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-66,-13,-66,-12.5</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-77,-16,-77,-13</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<intersection>-13 1</intersection></vsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-68.5,-21,-68.5,-14.5</points>
<intersection>-21 3</intersection>
<intersection>-17 1</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-71,-17,-68.5,-17</points>
<connection>
<GID>302</GID>
<name>OUT</name></connection>
<intersection>-68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-68.5,-14.5,-66,-14.5</points>
<connection>
<GID>303</GID>
<name>IN_1</name></connection>
<intersection>-68.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-68.5,-21,-66,-21</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<intersection>-68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-59.5,-16.5,-59.5,-13.5</points>
<intersection>-16.5 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-59.5,-16.5,-59,-16.5</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>-59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-60,-13.5,-59.5,-13.5</points>
<connection>
<GID>303</GID>
<name>OUT</name></connection>
<intersection>-59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-59.5,-22,-59.5,-18.5</points>
<intersection>-22 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-59.5,-18.5,-59,-18.5</points>
<connection>
<GID>305</GID>
<name>IN_1</name></connection>
<intersection>-59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-60,-22,-59.5,-22</points>
<connection>
<GID>304</GID>
<name>OUT</name></connection>
<intersection>-59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52.5,-18.5,-52.5,-16.5</points>
<intersection>-18.5 3</intersection>
<intersection>-17.5 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-52.5,-16.5,-52,-16.5</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<intersection>-52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-53,-17.5,-52.5,-17.5</points>
<connection>
<GID>305</GID>
<name>OUT</name></connection>
<intersection>-52.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-52.5,-18.5,-52,-18.5</points>
<connection>
<GID>306</GID>
<name>IN_1</name></connection>
<intersection>-52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-46,-17.5,-42.5,-17.5</points>
<connection>
<GID>306</GID>
<name>OUT</name></connection>
<intersection>-42.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-42.5,-18.5,-42.5,-16.5</points>
<connection>
<GID>307</GID>
<name>IN_1</name></connection>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>-17.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-36.5,-17.5,-27,-17.5</points>
<connection>
<GID>307</GID>
<name>OUT</name></connection>
<connection>
<GID>295</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>32.5081,-30.6493,101.436,-64.719</PageViewport>
<gate>
<ID>386</ID>
<type>AA_LABEL</type>
<position>54.5,-138.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>387</ID>
<type>AA_LABEL</type>
<position>60.5,-138.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>388</ID>
<type>AA_LABEL</type>
<position>63,-137</position>
<gparam>LABEL_TEXT __</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>389</ID>
<type>AA_LABEL</type>
<position>50,-137</position>
<gparam>LABEL_TEXT __</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>393</ID>
<type>BA_NAND2</type>
<position>48,-143.5</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>155 </input>
<output>
<ID>OUT</ID>158 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>394</ID>
<type>BA_NAND2</type>
<position>61,-143</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>156 </input>
<output>
<ID>OUT</ID>159 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>396</ID>
<type>BA_NAND2</type>
<position>72.5,-151.5</position>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_1</ID>156 </input>
<output>
<ID>OUT</ID>160 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>398</ID>
<type>BA_NAND2</type>
<position>73,-160</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>159 </input>
<output>
<ID>OUT</ID>161 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>400</ID>
<type>BA_NAND2</type>
<position>72.5,-167</position>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_1</ID>159 </input>
<output>
<ID>OUT</ID>157 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>401</ID>
<type>BA_NAND2</type>
<position>82.5,-155.5</position>
<input>
<ID>IN_0</ID>160 </input>
<input>
<ID>IN_1</ID>161 </input>
<output>
<ID>OUT</ID>167 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>402</ID>
<type>BA_NAND2</type>
<position>85,-167</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>157 </input>
<output>
<ID>OUT</ID>205 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>404</ID>
<type>GA_LED</type>
<position>94,-65.5</position>
<input>
<ID>N_in0</ID>166 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>406</ID>
<type>GA_LED</type>
<position>100,-120.5</position>
<input>
<ID>N_in0</ID>165 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>408</ID>
<type>GA_LED</type>
<position>104,-161</position>
<input>
<ID>N_in0</ID>167 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>410</ID>
<type>AA_LABEL</type>
<position>22.5,-43</position>
<gparam>LABEL_TEXT AOI</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>413</ID>
<type>AA_LABEL</type>
<position>158.5,-19.5</position>
<gparam>LABEL_TEXT Half Subtractor</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>414</ID>
<type>AA_TOGGLE</type>
<position>127.5,-27.5</position>
<output>
<ID>OUT_0</ID>168 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>415</ID>
<type>AA_TOGGLE</type>
<position>151,-27.5</position>
<output>
<ID>OUT_0</ID>169 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>416</ID>
<type>AA_AND2</type>
<position>166,-49.5</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>169 </input>
<output>
<ID>OUT</ID>172 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>417</ID>
<type>AA_AND2</type>
<position>166.5,-59.5</position>
<input>
<ID>IN_0</ID>168 </input>
<input>
<ID>IN_1</ID>171 </input>
<output>
<ID>OUT</ID>173 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>418</ID>
<type>AA_INVERTER</type>
<position>135.5,-35.5</position>
<input>
<ID>IN_0</ID>168 </input>
<output>
<ID>OUT_0</ID>170 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>419</ID>
<type>AA_INVERTER</type>
<position>157.5,-34.5</position>
<input>
<ID>IN_0</ID>169 </input>
<output>
<ID>OUT_0</ID>171 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>420</ID>
<type>GA_LED</type>
<position>198.5,-52.5</position>
<input>
<ID>N_in0</ID>174 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>421</ID>
<type>GA_LED</type>
<position>197.5,-64</position>
<input>
<ID>N_in0</ID>179 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>422</ID>
<type>AE_OR2</type>
<position>179.5,-52</position>
<input>
<ID>IN_0</ID>172 </input>
<input>
<ID>IN_1</ID>173 </input>
<output>
<ID>OUT</ID>174 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>423</ID>
<type>GA_LED</type>
<position>168.5,-79</position>
<input>
<ID>N_in1</ID>178 </input>
<input>
<ID>N_in2</ID>178 </input>
<input>
<ID>N_in3</ID>178 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>424</ID>
<type>GA_LED</type>
<position>168.5,-87.5</position>
<input>
<ID>N_in0</ID>177 </input>
<input>
<ID>N_in3</ID>177 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>425</ID>
<type>AI_XOR2</type>
<position>163,-79</position>
<input>
<ID>IN_0</ID>175 </input>
<input>
<ID>IN_1</ID>176 </input>
<output>
<ID>OUT</ID>178 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>426</ID>
<type>AA_TOGGLE</type>
<position>146.5,-77.5</position>
<output>
<ID>OUT_0</ID>175 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>427</ID>
<type>AA_TOGGLE</type>
<position>143.5,-80</position>
<output>
<ID>OUT_0</ID>176 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>428</ID>
<type>AA_AND2</type>
<position>165,-68</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>169 </input>
<output>
<ID>OUT</ID>179 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>429</ID>
<type>AA_AND2</type>
<position>162.5,-87.5</position>
<input>
<ID>IN_0</ID>180 </input>
<input>
<ID>IN_1</ID>176 </input>
<output>
<ID>OUT</ID>177 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>430</ID>
<type>AE_SMALL_INVERTER</type>
<position>154.5,-86.5</position>
<input>
<ID>IN_0</ID>175 </input>
<output>
<ID>OUT_0</ID>180 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>449</ID>
<type>AA_LABEL</type>
<position>140,-102</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>450</ID>
<type>AA_LABEL</type>
<position>146,-102</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>451</ID>
<type>AA_LABEL</type>
<position>148.5,-100.5</position>
<gparam>LABEL_TEXT __</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>452</ID>
<type>AA_LABEL</type>
<position>135.5,-100.5</position>
<gparam>LABEL_TEXT __</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>453</ID>
<type>BA_NAND2</type>
<position>133.5,-107</position>
<input>
<ID>IN_0</ID>187 </input>
<input>
<ID>IN_1</ID>187 </input>
<output>
<ID>OUT</ID>190 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>454</ID>
<type>BA_NAND2</type>
<position>146.5,-106.5</position>
<input>
<ID>IN_0</ID>188 </input>
<input>
<ID>IN_1</ID>188 </input>
<output>
<ID>OUT</ID>191 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>455</ID>
<type>BA_NAND2</type>
<position>158,-115</position>
<input>
<ID>IN_0</ID>190 </input>
<input>
<ID>IN_1</ID>188 </input>
<output>
<ID>OUT</ID>192 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>456</ID>
<type>BA_NAND2</type>
<position>158.5,-123.5</position>
<input>
<ID>IN_0</ID>187 </input>
<input>
<ID>IN_1</ID>191 </input>
<output>
<ID>OUT</ID>193 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>457</ID>
<type>BA_NAND2</type>
<position>158,-130.5</position>
<input>
<ID>IN_0</ID>190 </input>
<input>
<ID>IN_1</ID>188 </input>
<output>
<ID>OUT</ID>189 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>458</ID>
<type>BA_NAND2</type>
<position>168,-119</position>
<input>
<ID>IN_0</ID>192 </input>
<input>
<ID>IN_1</ID>193 </input>
<output>
<ID>OUT</ID>194 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>459</ID>
<type>BA_NAND2</type>
<position>170.5,-130.5</position>
<input>
<ID>IN_0</ID>189 </input>
<input>
<ID>IN_1</ID>189 </input>
<output>
<ID>OUT</ID>204 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>460</ID>
<type>GA_LED</type>
<position>189.5,-124.5</position>
<input>
<ID>N_in0</ID>194 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>461</ID>
<type>AA_LABEL</type>
<position>140.5,-96</position>
<gparam>LABEL_TEXT NAND IMPLEMENTATION</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>462</ID>
<type>AA_TOGGLE</type>
<position>127,-105</position>
<output>
<ID>OUT_0</ID>187 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>463</ID>
<type>AA_TOGGLE</type>
<position>140,-104.5</position>
<output>
<ID>OUT_0</ID>188 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>464</ID>
<type>AA_LABEL</type>
<position>127,-102</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>465</ID>
<type>AA_LABEL</type>
<position>133.5,-102</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>466</ID>
<type>GA_LED</type>
<position>184.5,-174</position>
<input>
<ID>N_in0</ID>202 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>467</ID>
<type>AA_LABEL</type>
<position>140.5,-140</position>
<gparam>LABEL_TEXT NOR IMPLEMENTATION</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>468</ID>
<type>AA_TOGGLE</type>
<position>124.5,-150</position>
<output>
<ID>OUT_0</ID>195 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>469</ID>
<type>AA_TOGGLE</type>
<position>137.5,-149.5</position>
<output>
<ID>OUT_0</ID>196 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>470</ID>
<type>AA_LABEL</type>
<position>124.5,-147</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>471</ID>
<type>AA_LABEL</type>
<position>131,-147</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>472</ID>
<type>AA_LABEL</type>
<position>137.5,-147</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>473</ID>
<type>AA_LABEL</type>
<position>143.5,-147</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>474</ID>
<type>AE_OR2</type>
<position>153.5,-158</position>
<input>
<ID>IN_0</ID>195 </input>
<input>
<ID>IN_1</ID>197 </input>
<output>
<ID>OUT</ID>199 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>475</ID>
<type>AE_OR2</type>
<position>154,-167</position>
<input>
<ID>IN_0</ID>198 </input>
<input>
<ID>IN_1</ID>196 </input>
<output>
<ID>OUT</ID>200 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>476</ID>
<type>AE_OR2</type>
<position>154,-176.5</position>
<input>
<ID>IN_0</ID>195 </input>
<input>
<ID>IN_1</ID>197 </input>
<output>
<ID>OUT</ID>203 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>477</ID>
<type>AE_OR2</type>
<position>170,-161.5</position>
<input>
<ID>IN_0</ID>199 </input>
<input>
<ID>IN_1</ID>200 </input>
<output>
<ID>OUT</ID>201 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>478</ID>
<type>AA_LABEL</type>
<position>146,-145.5</position>
<gparam>LABEL_TEXT __</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>479</ID>
<type>AA_LABEL</type>
<position>133,-145.5</position>
<gparam>LABEL_TEXT __</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>480</ID>
<type>BE_NOR2</type>
<position>131.5,-152</position>
<input>
<ID>IN_0</ID>195 </input>
<input>
<ID>IN_1</ID>195 </input>
<output>
<ID>OUT</ID>198 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>481</ID>
<type>BE_NOR2</type>
<position>144.5,-151.5</position>
<input>
<ID>IN_0</ID>196 </input>
<input>
<ID>IN_1</ID>196 </input>
<output>
<ID>OUT</ID>197 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>482</ID>
<type>BE_NOR2</type>
<position>181.5,-161.5</position>
<input>
<ID>IN_0</ID>201 </input>
<input>
<ID>IN_1</ID>201 </input>
<output>
<ID>OUT</ID>202 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>484</ID>
<type>GA_LED</type>
<position>176.5,-176.5</position>
<input>
<ID>N_in0</ID>203 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>486</ID>
<type>GA_LED</type>
<position>191,-130.5</position>
<input>
<ID>N_in0</ID>204 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>488</ID>
<type>GA_LED</type>
<position>104,-168.5</position>
<input>
<ID>N_in0</ID>205 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>490</ID>
<type>GA_LED</type>
<position>87,-123</position>
<input>
<ID>N_in0</ID>206 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>492</ID>
<type>GA_LED</type>
<position>99,-73.5</position>
<input>
<ID>N_in0</ID>207 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>310</ID>
<type>AA_LABEL</type>
<position>54,-17.5</position>
<gparam>LABEL_TEXT Half Adder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>314</ID>
<type>AI_XOR2</type>
<position>54.5,-29</position>
<input>
<ID>IN_0</ID>138 </input>
<input>
<ID>IN_1</ID>139 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>316</ID>
<type>AA_AND2</type>
<position>54,-36.5</position>
<input>
<ID>IN_0</ID>138 </input>
<input>
<ID>IN_1</ID>139 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>318</ID>
<type>AA_TOGGLE</type>
<position>40.5,-27</position>
<output>
<ID>OUT_0</ID>138 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>320</ID>
<type>AA_TOGGLE</type>
<position>40.5,-31</position>
<output>
<ID>OUT_0</ID>139 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>321</ID>
<type>AA_LABEL</type>
<position>63.5,-28.5</position>
<gparam>LABEL_TEXT Y = A.B + A.B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>322</ID>
<type>AA_LABEL</type>
<position>62,-27</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>323</ID>
<type>AA_LABEL</type>
<position>68,-27</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>324</ID>
<type>AA_LABEL</type>
<position>61,-36</position>
<gparam>LABEL_TEXT Y = A.B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>326</ID>
<type>AA_TOGGLE</type>
<position>41.5,-46</position>
<output>
<ID>OUT_0</ID>142 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>328</ID>
<type>AA_TOGGLE</type>
<position>54,-46.5</position>
<output>
<ID>OUT_0</ID>141 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>332</ID>
<type>AE_SMALL_INVERTER</type>
<position>47,-49</position>
<input>
<ID>IN_0</ID>142 </input>
<output>
<ID>OUT_0</ID>140 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>333</ID>
<type>AE_SMALL_INVERTER</type>
<position>60,-48.5</position>
<input>
<ID>IN_0</ID>141 </input>
<output>
<ID>OUT_0</ID>143 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>335</ID>
<type>AA_LABEL</type>
<position>41.5,-43</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>337</ID>
<type>AA_LABEL</type>
<position>48,-43</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>339</ID>
<type>AA_LABEL</type>
<position>50,-41.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>340</ID>
<type>AA_LABEL</type>
<position>54.5,-43</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>342</ID>
<type>AA_LABEL</type>
<position>63,-41.5</position>
<gparam>LABEL_TEXT __</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>343</ID>
<type>AA_LABEL</type>
<position>60.5,-43</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>344</ID>
<type>AA_AND2</type>
<position>71.5,-53.5</position>
<input>
<ID>IN_0</ID>140 </input>
<input>
<ID>IN_1</ID>141 </input>
<output>
<ID>OUT</ID>144 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>345</ID>
<type>AA_AND2</type>
<position>71.5,-63</position>
<input>
<ID>IN_0</ID>142 </input>
<input>
<ID>IN_1</ID>143 </input>
<output>
<ID>OUT</ID>145 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>347</ID>
<type>AE_OR2</type>
<position>85,-58</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>145 </input>
<output>
<ID>OUT</ID>166 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>349</ID>
<type>AA_AND2</type>
<position>71.5,-72</position>
<input>
<ID>IN_0</ID>142 </input>
<input>
<ID>IN_1</ID>141 </input>
<output>
<ID>OUT</ID>207 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>350</ID>
<type>AA_LABEL</type>
<position>94.5,-58</position>
<gparam>LABEL_TEXT Y = A.B + A.B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>351</ID>
<type>AA_LABEL</type>
<position>93,-56.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>352</ID>
<type>AA_LABEL</type>
<position>99,-56.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>353</ID>
<type>AA_LABEL</type>
<position>78,-71.5</position>
<gparam>LABEL_TEXT Y = A.B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>354</ID>
<type>AA_LABEL</type>
<position>79.5,-70</position>
<gparam>LABEL_TEXT ___</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>356</ID>
<type>AA_LABEL</type>
<position>56,-86.5</position>
<gparam>LABEL_TEXT NOR IMPLEMENTATION</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>357</ID>
<type>AA_TOGGLE</type>
<position>40,-96.5</position>
<output>
<ID>OUT_0</ID>146 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>358</ID>
<type>AA_TOGGLE</type>
<position>53,-96</position>
<output>
<ID>OUT_0</ID>147 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>361</ID>
<type>AA_LABEL</type>
<position>40,-93.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>362</ID>
<type>AA_LABEL</type>
<position>46.5,-93.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>363</ID>
<type>AA_LABEL</type>
<position>53,-93.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>364</ID>
<type>AA_LABEL</type>
<position>59,-93.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>366</ID>
<type>AE_OR2</type>
<position>69,-104.5</position>
<input>
<ID>IN_0</ID>146 </input>
<input>
<ID>IN_1</ID>148 </input>
<output>
<ID>OUT</ID>150 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>368</ID>
<type>AE_OR2</type>
<position>69.5,-113.5</position>
<input>
<ID>IN_0</ID>149 </input>
<input>
<ID>IN_1</ID>147 </input>
<output>
<ID>OUT</ID>151 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>370</ID>
<type>AE_OR2</type>
<position>69.5,-123</position>
<input>
<ID>IN_0</ID>149 </input>
<input>
<ID>IN_1</ID>148 </input>
<output>
<ID>OUT</ID>206 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>372</ID>
<type>AE_OR2</type>
<position>85.5,-108</position>
<input>
<ID>IN_0</ID>150 </input>
<input>
<ID>IN_1</ID>151 </input>
<output>
<ID>OUT</ID>152 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>375</ID>
<type>AA_LABEL</type>
<position>61.5,-92</position>
<gparam>LABEL_TEXT __</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>376</ID>
<type>AA_LABEL</type>
<position>48.5,-92</position>
<gparam>LABEL_TEXT __</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>378</ID>
<type>BE_NOR2</type>
<position>47,-98.5</position>
<input>
<ID>IN_0</ID>146 </input>
<input>
<ID>IN_1</ID>146 </input>
<output>
<ID>OUT</ID>149 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>379</ID>
<type>BE_NOR2</type>
<position>60,-98</position>
<input>
<ID>IN_0</ID>147 </input>
<input>
<ID>IN_1</ID>147 </input>
<output>
<ID>OUT</ID>148 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>380</ID>
<type>BE_NOR2</type>
<position>97,-108</position>
<input>
<ID>IN_0</ID>152 </input>
<input>
<ID>IN_1</ID>152 </input>
<output>
<ID>OUT</ID>165 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>381</ID>
<type>AA_LABEL</type>
<position>55,-132.5</position>
<gparam>LABEL_TEXT NAND IMPLEMENTATION</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>382</ID>
<type>AA_TOGGLE</type>
<position>41.5,-141.5</position>
<output>
<ID>OUT_0</ID>155 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>383</ID>
<type>AA_TOGGLE</type>
<position>54.5,-141</position>
<output>
<ID>OUT_0</ID>156 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>384</ID>
<type>AA_LABEL</type>
<position>41.5,-138.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>385</ID>
<type>AA_LABEL</type>
<position>48,-138.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,-123.5,163,-120</points>
<intersection>-123.5 1</intersection>
<intersection>-120 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161.5,-123.5,163,-123.5</points>
<connection>
<GID>456</GID>
<name>OUT</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>163,-120,165,-120</points>
<connection>
<GID>458</GID>
<name>IN_1</name></connection>
<intersection>163 0</intersection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179.5,-124.5,179.5,-119</points>
<intersection>-124.5 2</intersection>
<intersection>-119 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>171,-119,179.5,-119</points>
<connection>
<GID>458</GID>
<name>OUT</name></connection>
<intersection>179.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>179.5,-124.5,188.5,-124.5</points>
<connection>
<GID>460</GID>
<name>N_in0</name></connection>
<intersection>179.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-175.5,124.5,-152</points>
<connection>
<GID>468</GID>
<name>OUT_0</name></connection>
<intersection>-175.5 7</intersection>
<intersection>-157 1</intersection>
<intersection>-152 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124.5,-157,150.5,-157</points>
<connection>
<GID>474</GID>
<name>IN_0</name></connection>
<intersection>124.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124.5,-152,128,-152</points>
<intersection>124.5 0</intersection>
<intersection>128 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>128,-153,128,-151</points>
<intersection>-153 5</intersection>
<intersection>-152 2</intersection>
<intersection>-151 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>128,-151,128.5,-151</points>
<connection>
<GID>480</GID>
<name>IN_0</name></connection>
<intersection>128 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>128,-153,128.5,-153</points>
<connection>
<GID>480</GID>
<name>IN_1</name></connection>
<intersection>128 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>124.5,-175.5,151,-175.5</points>
<connection>
<GID>476</GID>
<name>IN_0</name></connection>
<intersection>124.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>140.5,-152.5,140.5,-150.5</points>
<intersection>-152.5 13</intersection>
<intersection>-151.5 5</intersection>
<intersection>-150.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>140.5,-150.5,141.5,-150.5</points>
<connection>
<GID>481</GID>
<name>IN_0</name></connection>
<intersection>140.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>137.5,-151.5,140.5,-151.5</points>
<intersection>137.5 8</intersection>
<intersection>140.5 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>137.5,-168,137.5,-151.5</points>
<connection>
<GID>469</GID>
<name>OUT_0</name></connection>
<intersection>-168 11</intersection>
<intersection>-151.5 5</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>137.5,-168,151,-168</points>
<connection>
<GID>475</GID>
<name>IN_1</name></connection>
<intersection>137.5 8</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>140.5,-152.5,141.5,-152.5</points>
<connection>
<GID>481</GID>
<name>IN_1</name></connection>
<intersection>140.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149,-177.5,149,-151.5</points>
<intersection>-177.5 4</intersection>
<intersection>-159 1</intersection>
<intersection>-151.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>149,-159,150.5,-159</points>
<connection>
<GID>474</GID>
<name>IN_1</name></connection>
<intersection>149 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>147.5,-151.5,149,-151.5</points>
<connection>
<GID>481</GID>
<name>OUT</name></connection>
<intersection>149 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>149,-177.5,151,-177.5</points>
<connection>
<GID>476</GID>
<name>IN_1</name></connection>
<intersection>149 0</intersection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134.5,-166,134.5,-152</points>
<connection>
<GID>480</GID>
<name>OUT</name></connection>
<intersection>-166 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>134.5,-166,151,-166</points>
<connection>
<GID>475</GID>
<name>IN_0</name></connection>
<intersection>134.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161.5,-160.5,161.5,-158</points>
<intersection>-160.5 2</intersection>
<intersection>-158 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156.5,-158,161.5,-158</points>
<connection>
<GID>474</GID>
<name>OUT</name></connection>
<intersection>161.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>161.5,-160.5,167,-160.5</points>
<connection>
<GID>477</GID>
<name>IN_0</name></connection>
<intersection>161.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-167,162,-162.5</points>
<intersection>-167 1</intersection>
<intersection>-162.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157,-167,162,-167</points>
<connection>
<GID>475</GID>
<name>OUT</name></connection>
<intersection>162 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162,-162.5,167,-162.5</points>
<connection>
<GID>477</GID>
<name>IN_1</name></connection>
<intersection>162 0</intersection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>177.5,-162.5,177.5,-160.5</points>
<intersection>-162.5 13</intersection>
<intersection>-161.5 14</intersection>
<intersection>-160.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>177.5,-160.5,178.5,-160.5</points>
<connection>
<GID>482</GID>
<name>IN_0</name></connection>
<intersection>177.5 3</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>177.5,-162.5,178.5,-162.5</points>
<connection>
<GID>482</GID>
<name>IN_1</name></connection>
<intersection>177.5 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>173,-161.5,177.5,-161.5</points>
<connection>
<GID>477</GID>
<name>OUT</name></connection>
<intersection>177.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,-174,184,-161.5</points>
<intersection>-174 2</intersection>
<intersection>-161.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,-161.5,184.5,-161.5</points>
<connection>
<GID>482</GID>
<name>OUT</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>183.5,-174,184,-174</points>
<connection>
<GID>466</GID>
<name>N_in0</name></connection>
<intersection>184 0</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,-176.5,175.5,-176.5</points>
<connection>
<GID>476</GID>
<name>OUT</name></connection>
<connection>
<GID>484</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>173.5,-130.5,190,-130.5</points>
<connection>
<GID>459</GID>
<name>OUT</name></connection>
<connection>
<GID>486</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-168.5,95.5,-167</points>
<intersection>-168.5 2</intersection>
<intersection>-167 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88,-167,95.5,-167</points>
<connection>
<GID>402</GID>
<name>OUT</name></connection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95.5,-168.5,103,-168.5</points>
<connection>
<GID>488</GID>
<name>N_in0</name></connection>
<intersection>95.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72.5,-123,86,-123</points>
<connection>
<GID>370</GID>
<name>OUT</name></connection>
<connection>
<GID>490</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-73.5,86,-72</points>
<intersection>-73.5 2</intersection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-72,86,-72</points>
<connection>
<GID>349</GID>
<name>OUT</name></connection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86,-73.5,98,-73.5</points>
<connection>
<GID>492</GID>
<name>N_in0</name></connection>
<intersection>86 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42.5,-27,51.5,-27</points>
<connection>
<GID>318</GID>
<name>OUT_0</name></connection>
<intersection>44.5 6</intersection>
<intersection>51.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>51.5,-28,51.5,-27</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<intersection>-27 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>44.5,-35.5,44.5,-27</points>
<intersection>-35.5 7</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>44.5,-35.5,51,-35.5</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>44.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42.5,-31,51.5,-31</points>
<connection>
<GID>320</GID>
<name>OUT_0</name></connection>
<intersection>46.5 5</intersection>
<intersection>51.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>51.5,-31,51.5,-30</points>
<connection>
<GID>314</GID>
<name>IN_1</name></connection>
<intersection>-31 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>46.5,-37.5,46.5,-31</points>
<intersection>-37.5 6</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>46.5,-37.5,51,-37.5</points>
<connection>
<GID>316</GID>
<name>IN_1</name></connection>
<intersection>46.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-52.5,47,-51</points>
<connection>
<GID>332</GID>
<name>OUT_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-52.5,68.5,-52.5</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-73,54,-46.5</points>
<connection>
<GID>328</GID>
<name>OUT_0</name></connection>
<intersection>-73 3</intersection>
<intersection>-54.5 1</intersection>
<intersection>-46.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-54.5,68.5,-54.5</points>
<connection>
<GID>344</GID>
<name>IN_1</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>54,-73,68.5,-73</points>
<connection>
<GID>349</GID>
<name>IN_1</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>54,-46.5,60,-46.5</points>
<connection>
<GID>333</GID>
<name>IN_0</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-71,41.5,-47.5</points>
<connection>
<GID>326</GID>
<name>OUT_0</name></connection>
<intersection>-71 3</intersection>
<intersection>-62 1</intersection>
<intersection>-47.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-62,68.5,-62</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>41.5,-71,68.5,-71</points>
<connection>
<GID>349</GID>
<name>IN_0</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>41.5,-47.5,47,-47.5</points>
<intersection>41.5 0</intersection>
<intersection>47 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>47,-47.5,47,-47</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<intersection>-47.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-64,60,-50.5</points>
<connection>
<GID>333</GID>
<name>OUT_0</name></connection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60,-64,68.5,-64</points>
<connection>
<GID>345</GID>
<name>IN_1</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-57,78,-53.5</points>
<intersection>-57 2</intersection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-53.5,78,-53.5</points>
<connection>
<GID>344</GID>
<name>OUT</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78,-57,82,-57</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-63,78,-59</points>
<intersection>-63 1</intersection>
<intersection>-59 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-63,78,-63</points>
<connection>
<GID>345</GID>
<name>OUT</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78,-59,82,-59</points>
<connection>
<GID>347</GID>
<name>IN_1</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-103.5,40,-98.5</points>
<connection>
<GID>357</GID>
<name>OUT_0</name></connection>
<intersection>-103.5 1</intersection>
<intersection>-98.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-103.5,66,-103.5</points>
<connection>
<GID>366</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40,-98.5,43.5,-98.5</points>
<intersection>40 0</intersection>
<intersection>43.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>43.5,-99.5,43.5,-97.5</points>
<intersection>-99.5 5</intersection>
<intersection>-98.5 2</intersection>
<intersection>-97.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>43.5,-97.5,44,-97.5</points>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<intersection>43.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>43.5,-99.5,44,-99.5</points>
<connection>
<GID>378</GID>
<name>IN_1</name></connection>
<intersection>43.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>56,-99,56,-97</points>
<intersection>-99 13</intersection>
<intersection>-98 5</intersection>
<intersection>-97 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>56,-97,57,-97</points>
<connection>
<GID>379</GID>
<name>IN_0</name></connection>
<intersection>56 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>53,-98,56,-98</points>
<intersection>53 8</intersection>
<intersection>56 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>53,-114.5,53,-98</points>
<connection>
<GID>358</GID>
<name>OUT_0</name></connection>
<intersection>-114.5 11</intersection>
<intersection>-98 5</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>53,-114.5,66.5,-114.5</points>
<connection>
<GID>368</GID>
<name>IN_1</name></connection>
<intersection>53 8</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>56,-99,57,-99</points>
<connection>
<GID>379</GID>
<name>IN_1</name></connection>
<intersection>56 3</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-124,64.5,-98</points>
<intersection>-124 4</intersection>
<intersection>-105.5 1</intersection>
<intersection>-98 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64.5,-105.5,66,-105.5</points>
<connection>
<GID>366</GID>
<name>IN_1</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63,-98,64.5,-98</points>
<connection>
<GID>379</GID>
<name>OUT</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>64.5,-124,66.5,-124</points>
<connection>
<GID>370</GID>
<name>IN_1</name></connection>
<intersection>64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-122,50,-98.5</points>
<connection>
<GID>378</GID>
<name>OUT</name></connection>
<intersection>-122 4</intersection>
<intersection>-112.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>50,-112.5,66.5,-112.5</points>
<connection>
<GID>368</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>50,-122,66.5,-122</points>
<connection>
<GID>370</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-107,77,-104.5</points>
<intersection>-107 2</intersection>
<intersection>-104.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-104.5,77,-104.5</points>
<connection>
<GID>366</GID>
<name>OUT</name></connection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-107,82.5,-107</points>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-113.5,77.5,-109</points>
<intersection>-113.5 1</intersection>
<intersection>-109 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-113.5,77.5,-113.5</points>
<connection>
<GID>368</GID>
<name>OUT</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77.5,-109,82.5,-109</points>
<connection>
<GID>372</GID>
<name>IN_1</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>93,-109,93,-107</points>
<intersection>-109 13</intersection>
<intersection>-108 14</intersection>
<intersection>-107 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>93,-107,94,-107</points>
<connection>
<GID>380</GID>
<name>IN_0</name></connection>
<intersection>93 3</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>93,-109,94,-109</points>
<connection>
<GID>380</GID>
<name>IN_1</name></connection>
<intersection>93 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>88.5,-108,93,-108</points>
<connection>
<GID>372</GID>
<name>OUT</name></connection>
<intersection>93 3</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-159,41.5,-143.5</points>
<connection>
<GID>382</GID>
<name>OUT_0</name></connection>
<intersection>-159 8</intersection>
<intersection>-143.5 9</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>41.5,-159,70,-159</points>
<connection>
<GID>398</GID>
<name>IN_0</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>41.5,-143.5,45,-143.5</points>
<intersection>41.5 0</intersection>
<intersection>45 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>45,-144.5,45,-142.5</points>
<connection>
<GID>393</GID>
<name>IN_0</name></connection>
<connection>
<GID>393</GID>
<name>IN_1</name></connection>
<intersection>-143.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-152.5,54.5,-143</points>
<connection>
<GID>383</GID>
<name>OUT_0</name></connection>
<intersection>-152.5 4</intersection>
<intersection>-143 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>54.5,-152.5,69.5,-152.5</points>
<connection>
<GID>396</GID>
<name>IN_1</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>54.5,-143,58,-143</points>
<intersection>54.5 0</intersection>
<intersection>58 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>58,-144,58,-142</points>
<connection>
<GID>394</GID>
<name>IN_1</name></connection>
<connection>
<GID>394</GID>
<name>IN_0</name></connection>
<intersection>-143 5</intersection></vsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-168,82,-166</points>
<connection>
<GID>402</GID>
<name>IN_1</name></connection>
<connection>
<GID>402</GID>
<name>IN_0</name></connection>
<intersection>-167 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75.5,-167,82,-167</points>
<connection>
<GID>400</GID>
<name>OUT</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-166,52,-143.5</points>
<intersection>-166 4</intersection>
<intersection>-150.5 2</intersection>
<intersection>-143.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-143.5,52,-143.5</points>
<connection>
<GID>393</GID>
<name>OUT</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,-150.5,69.5,-150.5</points>
<connection>
<GID>396</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>52,-166,69.5,-166</points>
<connection>
<GID>400</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-168,67,-143</points>
<intersection>-168 4</intersection>
<intersection>-161 2</intersection>
<intersection>-143 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,-143,67,-143</points>
<connection>
<GID>394</GID>
<name>OUT</name></connection>
<intersection>67 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>67,-161,70,-161</points>
<connection>
<GID>398</GID>
<name>IN_1</name></connection>
<intersection>67 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>67,-168,69.5,-168</points>
<connection>
<GID>400</GID>
<name>IN_1</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-154.5,77.5,-151.5</points>
<intersection>-154.5 2</intersection>
<intersection>-151.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75.5,-151.5,77.5,-151.5</points>
<connection>
<GID>396</GID>
<name>OUT</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77.5,-154.5,79.5,-154.5</points>
<connection>
<GID>401</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-160,77.5,-156.5</points>
<intersection>-160 1</intersection>
<intersection>-156.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-160,77.5,-160</points>
<connection>
<GID>398</GID>
<name>OUT</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77.5,-156.5,79.5,-156.5</points>
<connection>
<GID>401</GID>
<name>IN_1</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-120.5,99.5,-108</points>
<intersection>-120.5 2</intersection>
<intersection>-108 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99.5,-108,100,-108</points>
<connection>
<GID>380</GID>
<name>OUT</name></connection>
<intersection>99.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-120.5,99.5,-120.5</points>
<connection>
<GID>406</GID>
<name>N_in0</name></connection>
<intersection>99.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-65.5,90.5,-58</points>
<intersection>-65.5 2</intersection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88,-58,90.5,-58</points>
<connection>
<GID>347</GID>
<name>OUT</name></connection>
<intersection>90.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-65.5,93,-65.5</points>
<connection>
<GID>404</GID>
<name>N_in0</name></connection>
<intersection>90.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94,-161,94,-155.5</points>
<intersection>-161 2</intersection>
<intersection>-155.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-155.5,94,-155.5</points>
<connection>
<GID>401</GID>
<name>OUT</name></connection>
<intersection>94 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94,-161,103,-161</points>
<connection>
<GID>408</GID>
<name>N_in0</name></connection>
<intersection>94 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,-58.5,127.5,-29.5</points>
<connection>
<GID>414</GID>
<name>OUT_0</name></connection>
<intersection>-58.5 3</intersection>
<intersection>-32.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>127.5,-58.5,163.5,-58.5</points>
<connection>
<GID>417</GID>
<name>IN_0</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>127.5,-32.5,135.5,-32.5</points>
<connection>
<GID>418</GID>
<name>IN_0</name></connection>
<intersection>127.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-50.5,151,-29.5</points>
<connection>
<GID>415</GID>
<name>OUT_0</name></connection>
<intersection>-50.5 2</intersection>
<intersection>-31.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>151,-50.5,163,-50.5</points>
<connection>
<GID>416</GID>
<name>IN_1</name></connection>
<intersection>151 0</intersection>
<intersection>151.5 5</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>151,-31.5,157.5,-31.5</points>
<connection>
<GID>419</GID>
<name>IN_0</name></connection>
<intersection>151 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>151.5,-69,151.5,-50.5</points>
<intersection>-69 6</intersection>
<intersection>-50.5 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>151.5,-69,162,-69</points>
<connection>
<GID>428</GID>
<name>IN_1</name></connection>
<intersection>151.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-48.5,135.5,-38.5</points>
<connection>
<GID>418</GID>
<name>OUT_0</name></connection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-48.5,163,-48.5</points>
<connection>
<GID>416</GID>
<name>IN_0</name></connection>
<intersection>135 2</intersection>
<intersection>135.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>135,-67,135,-48.5</points>
<intersection>-67 3</intersection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>135,-67,162,-67</points>
<connection>
<GID>428</GID>
<name>IN_0</name></connection>
<intersection>135 2</intersection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157.5,-60.5,157.5,-37.5</points>
<connection>
<GID>419</GID>
<name>OUT_0</name></connection>
<intersection>-60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,-60.5,163.5,-60.5</points>
<connection>
<GID>417</GID>
<name>IN_1</name></connection>
<intersection>157.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172.5,-51,172.5,-49.5</points>
<intersection>-51 1</intersection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172.5,-51,176.5,-51</points>
<connection>
<GID>422</GID>
<name>IN_0</name></connection>
<intersection>172.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>169,-49.5,172.5,-49.5</points>
<connection>
<GID>416</GID>
<name>OUT</name></connection>
<intersection>172.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173,-59.5,173,-53</points>
<intersection>-59.5 2</intersection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>173,-53,176.5,-53</points>
<connection>
<GID>422</GID>
<name>IN_1</name></connection>
<intersection>173 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>169.5,-59.5,173,-59.5</points>
<connection>
<GID>417</GID>
<name>OUT</name></connection>
<intersection>173 0</intersection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190,-52.5,190,-52</points>
<intersection>-52.5 1</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190,-52.5,197.5,-52.5</points>
<connection>
<GID>420</GID>
<name>N_in0</name></connection>
<intersection>190 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>182.5,-52,190,-52</points>
<connection>
<GID>422</GID>
<name>OUT</name></connection>
<intersection>190 0</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>148.5,-78,160,-78</points>
<connection>
<GID>425</GID>
<name>IN_0</name></connection>
<intersection>148.5 10</intersection>
<intersection>152.5 11</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>148.5,-78,148.5,-77.5</points>
<connection>
<GID>426</GID>
<name>OUT_0</name></connection>
<intersection>-78 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>152.5,-86.5,152.5,-78</points>
<connection>
<GID>430</GID>
<name>IN_0</name></connection>
<intersection>-78 1</intersection></vsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>145.5,-79.5,147,-79.5</points>
<intersection>145.5 7</intersection>
<intersection>147 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>147,-88.5,147,-79.5</points>
<intersection>-88.5 8</intersection>
<intersection>-80 9</intersection>
<intersection>-79.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>145.5,-80,145.5,-79.5</points>
<connection>
<GID>427</GID>
<name>OUT_0</name></connection>
<intersection>-79.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>147,-88.5,159.5,-88.5</points>
<connection>
<GID>429</GID>
<name>IN_1</name></connection>
<intersection>147 6</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>147,-80,160,-80</points>
<connection>
<GID>425</GID>
<name>IN_1</name></connection>
<intersection>147 6</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165.5,-87.5,168.5,-87.5</points>
<connection>
<GID>424</GID>
<name>N_in0</name></connection>
<connection>
<GID>429</GID>
<name>OUT</name></connection>
<intersection>168.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>168.5,-87.5,168.5,-86.5</points>
<connection>
<GID>424</GID>
<name>N_in3</name></connection>
<intersection>-87.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168.5,-80,168.5,-78</points>
<connection>
<GID>423</GID>
<name>N_in3</name></connection>
<connection>
<GID>423</GID>
<name>N_in2</name></connection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166,-79,169.5,-79</points>
<connection>
<GID>423</GID>
<name>N_in1</name></connection>
<connection>
<GID>425</GID>
<name>OUT</name></connection>
<intersection>168.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,-68,182,-64</points>
<intersection>-68 2</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>182,-64,196.5,-64</points>
<connection>
<GID>421</GID>
<name>N_in0</name></connection>
<intersection>182 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>168,-68,182,-68</points>
<connection>
<GID>428</GID>
<name>OUT</name></connection>
<intersection>182 0</intersection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,-86.5,159.5,-86.5</points>
<connection>
<GID>429</GID>
<name>IN_0</name></connection>
<connection>
<GID>430</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,-122.5,127,-107</points>
<connection>
<GID>462</GID>
<name>OUT_0</name></connection>
<intersection>-122.5 8</intersection>
<intersection>-107 9</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>127,-122.5,155.5,-122.5</points>
<connection>
<GID>456</GID>
<name>IN_0</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>127,-107,130.5,-107</points>
<intersection>127 0</intersection>
<intersection>130.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>130.5,-108,130.5,-106</points>
<connection>
<GID>453</GID>
<name>IN_1</name></connection>
<connection>
<GID>453</GID>
<name>IN_0</name></connection>
<intersection>-107 9</intersection></vsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,-131.5,140,-106.5</points>
<connection>
<GID>463</GID>
<name>OUT_0</name></connection>
<intersection>-131.5 12</intersection>
<intersection>-116 4</intersection>
<intersection>-106.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>140,-116,155,-116</points>
<connection>
<GID>455</GID>
<name>IN_1</name></connection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>140,-106.5,143.5,-106.5</points>
<intersection>140 0</intersection>
<intersection>143.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>143.5,-107.5,143.5,-105.5</points>
<connection>
<GID>454</GID>
<name>IN_1</name></connection>
<connection>
<GID>454</GID>
<name>IN_0</name></connection>
<intersection>-106.5 5</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>140,-131.5,155,-131.5</points>
<connection>
<GID>457</GID>
<name>IN_1</name></connection>
<intersection>140 0</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167.5,-131.5,167.5,-129.5</points>
<connection>
<GID>459</GID>
<name>IN_1</name></connection>
<connection>
<GID>459</GID>
<name>IN_0</name></connection>
<intersection>-130.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>161,-130.5,167.5,-130.5</points>
<connection>
<GID>457</GID>
<name>OUT</name></connection>
<intersection>167.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137.5,-129.5,137.5,-107</points>
<intersection>-129.5 4</intersection>
<intersection>-114 2</intersection>
<intersection>-107 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136.5,-107,137.5,-107</points>
<connection>
<GID>453</GID>
<name>OUT</name></connection>
<intersection>137.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>137.5,-114,155,-114</points>
<connection>
<GID>455</GID>
<name>IN_0</name></connection>
<intersection>137.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>137.5,-129.5,155,-129.5</points>
<connection>
<GID>457</GID>
<name>IN_0</name></connection>
<intersection>137.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152.5,-124.5,152.5,-106.5</points>
<intersection>-124.5 2</intersection>
<intersection>-106.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>149.5,-106.5,152.5,-106.5</points>
<connection>
<GID>454</GID>
<name>OUT</name></connection>
<intersection>152.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>152.5,-124.5,155.5,-124.5</points>
<connection>
<GID>456</GID>
<name>IN_1</name></connection>
<intersection>152.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,-118,163,-115</points>
<intersection>-118 2</intersection>
<intersection>-115 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161,-115,163,-115</points>
<connection>
<GID>455</GID>
<name>OUT</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>163,-118,165,-118</points>
<connection>
<GID>458</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>-35.6,-29.0372,182,-136.593</PageViewport>
<gate>
<ID>494</ID>
<type>AA_LABEL</type>
<position>39.5,-17.5</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>495</ID>
<type>AA_LABEL</type>
<position>186.5,-16</position>
<gparam>LABEL_TEXT Full Substractor</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>497</ID>
<type>AA_LABEL</type>
<position>37,-30.5</position>
<gparam>LABEL_TEXT AOI</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>507</ID>
<type>AA_TOGGLE</type>
<position>27.5,-38.5</position>
<output>
<ID>OUT_0</ID>220 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>508</ID>
<type>AA_TOGGLE</type>
<position>40,-39</position>
<output>
<ID>OUT_0</ID>209 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>509</ID>
<type>AE_SMALL_INVERTER</type>
<position>33,-42</position>
<input>
<ID>IN_0</ID>220 </input>
<output>
<ID>OUT_0</ID>217 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>510</ID>
<type>AE_SMALL_INVERTER</type>
<position>46.5,-42.5</position>
<input>
<ID>IN_0</ID>209 </input>
<output>
<ID>OUT_0</ID>218 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>511</ID>
<type>AA_LABEL</type>
<position>27.5,-35.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>512</ID>
<type>AA_LABEL</type>
<position>34,-35.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>513</ID>
<type>AA_LABEL</type>
<position>36,-34</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>514</ID>
<type>AA_LABEL</type>
<position>40.5,-35.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>515</ID>
<type>AA_LABEL</type>
<position>49,-34</position>
<gparam>LABEL_TEXT __</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>516</ID>
<type>AA_LABEL</type>
<position>46.5,-35.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>517</ID>
<type>AA_TOGGLE</type>
<position>55,-39</position>
<output>
<ID>OUT_0</ID>211 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>518</ID>
<type>AE_SMALL_INVERTER</type>
<position>62.5,-41.5</position>
<input>
<ID>IN_0</ID>211 </input>
<output>
<ID>OUT_0</ID>219 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>519</ID>
<type>AA_LABEL</type>
<position>55.5,-35.5</position>
<gparam>LABEL_TEXT Input Cin</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>520</ID>
<type>AA_LABEL</type>
<position>65.5,-36.5</position>
<gparam>LABEL_TEXT ____</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>521</ID>
<type>AA_LABEL</type>
<position>63,-38</position>
<gparam>LABEL_TEXT Input Cin</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>523</ID>
<type>AA_AND3</type>
<position>75,-48</position>
<input>
<ID>IN_0</ID>217 </input>
<input>
<ID>IN_1</ID>218 </input>
<input>
<ID>IN_2</ID>211 </input>
<output>
<ID>OUT</ID>221 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>525</ID>
<type>AA_AND3</type>
<position>75,-61.5</position>
<input>
<ID>IN_0</ID>217 </input>
<input>
<ID>IN_1</ID>209 </input>
<input>
<ID>IN_2</ID>219 </input>
<output>
<ID>OUT</ID>222 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>527</ID>
<type>AA_AND3</type>
<position>75,-72.5</position>
<input>
<ID>IN_0</ID>220 </input>
<input>
<ID>IN_1</ID>218 </input>
<input>
<ID>IN_2</ID>219 </input>
<output>
<ID>OUT</ID>223 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>529</ID>
<type>AA_AND3</type>
<position>75,-83</position>
<input>
<ID>IN_0</ID>220 </input>
<input>
<ID>IN_1</ID>209 </input>
<input>
<ID>IN_2</ID>211 </input>
<output>
<ID>OUT</ID>224 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>533</ID>
<type>GA_LED</type>
<position>107.5,-59</position>
<input>
<ID>N_in0</ID>225 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>535</ID>
<type>AE_OR4</type>
<position>94,-61</position>
<input>
<ID>IN_0</ID>221 </input>
<input>
<ID>IN_1</ID>222 </input>
<input>
<ID>IN_2</ID>223 </input>
<input>
<ID>IN_3</ID>224 </input>
<output>
<ID>OUT</ID>225 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>536</ID>
<type>AA_AND3</type>
<position>74.5,-95</position>
<input>
<ID>IN_0</ID>217 </input>
<input>
<ID>IN_1</ID>209 </input>
<input>
<ID>IN_2</ID>211 </input>
<output>
<ID>OUT</ID>227 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>537</ID>
<type>AA_AND3</type>
<position>75,-107.5</position>
<input>
<ID>IN_0</ID>220 </input>
<input>
<ID>IN_1</ID>218 </input>
<input>
<ID>IN_2</ID>211 </input>
<output>
<ID>OUT</ID>228 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>538</ID>
<type>AA_AND3</type>
<position>75.5,-119</position>
<input>
<ID>IN_0</ID>220 </input>
<input>
<ID>IN_1</ID>209 </input>
<input>
<ID>IN_2</ID>219 </input>
<output>
<ID>OUT</ID>229 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>539</ID>
<type>AA_AND3</type>
<position>75.5,-131.5</position>
<input>
<ID>IN_0</ID>220 </input>
<input>
<ID>IN_1</ID>209 </input>
<input>
<ID>IN_2</ID>211 </input>
<output>
<ID>OUT</ID>230 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>543</ID>
<type>GA_LED</type>
<position>110.5,-102</position>
<input>
<ID>N_in0</ID>226 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>544</ID>
<type>AE_OR4</type>
<position>97,-104</position>
<input>
<ID>IN_0</ID>227 </input>
<input>
<ID>IN_1</ID>228 </input>
<input>
<ID>IN_2</ID>229 </input>
<input>
<ID>IN_3</ID>230 </input>
<output>
<ID>OUT</ID>226 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<wire>
<ID>209</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>40,-41,46.5,-41</points>
<connection>
<GID>508</GID>
<name>OUT_0</name></connection>
<intersection>40 6</intersection>
<intersection>46.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>46.5,-41,46.5,-40.5</points>
<connection>
<GID>510</GID>
<name>IN_0</name></connection>
<intersection>-41 4</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>40,-131.5,40,-41</points>
<intersection>-131.5 17</intersection>
<intersection>-119 15</intersection>
<intersection>-95 13</intersection>
<intersection>-83 11</intersection>
<intersection>-61.5 7</intersection>
<intersection>-41 4</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>40,-61.5,72,-61.5</points>
<connection>
<GID>525</GID>
<name>IN_1</name></connection>
<intersection>40 6</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>40,-83,72,-83</points>
<connection>
<GID>529</GID>
<name>IN_1</name></connection>
<intersection>40 6</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>40,-95,71.5,-95</points>
<connection>
<GID>536</GID>
<name>IN_1</name></connection>
<intersection>40 6</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>40,-119,72.5,-119</points>
<connection>
<GID>538</GID>
<name>IN_1</name></connection>
<intersection>40 6</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>40,-131.5,72.5,-131.5</points>
<connection>
<GID>539</GID>
<name>IN_1</name></connection>
<intersection>40 6</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>7</ID>
<points>55,-133.5,55,-39.5</points>
<connection>
<GID>517</GID>
<name>OUT_0</name></connection>
<intersection>-133.5 18</intersection>
<intersection>-109.5 16</intersection>
<intersection>-97 14</intersection>
<intersection>-85 11</intersection>
<intersection>-50 12</intersection>
<intersection>-39.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>55,-39.5,62.5,-39.5</points>
<connection>
<GID>518</GID>
<name>IN_0</name></connection>
<intersection>55 7</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>55,-85,72,-85</points>
<connection>
<GID>529</GID>
<name>IN_2</name></connection>
<intersection>55 7</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>55,-50,72,-50</points>
<connection>
<GID>523</GID>
<name>IN_2</name></connection>
<intersection>55 7</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>55,-97,71.5,-97</points>
<connection>
<GID>536</GID>
<name>IN_2</name></connection>
<intersection>55 7</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>55,-109.5,72,-109.5</points>
<connection>
<GID>537</GID>
<name>IN_2</name></connection>
<intersection>55 7</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>55,-133.5,72.5,-133.5</points>
<connection>
<GID>539</GID>
<name>IN_2</name></connection>
<intersection>55 7</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-93,33,-44</points>
<connection>
<GID>509</GID>
<name>OUT_0</name></connection>
<intersection>-93 5</intersection>
<intersection>-59.5 3</intersection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-46,72,-46</points>
<connection>
<GID>523</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33,-59.5,72,-59.5</points>
<connection>
<GID>525</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>33,-93,71.5,-93</points>
<connection>
<GID>536</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-107.5,46.5,-44.5</points>
<connection>
<GID>510</GID>
<name>OUT_0</name></connection>
<intersection>-107.5 5</intersection>
<intersection>-72.5 3</intersection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-48,72,-48</points>
<connection>
<GID>523</GID>
<name>IN_1</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>46.5,-72.5,72,-72.5</points>
<connection>
<GID>527</GID>
<name>IN_1</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>46.5,-107.5,72,-107.5</points>
<connection>
<GID>537</GID>
<name>IN_1</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-121,62.5,-43.5</points>
<connection>
<GID>518</GID>
<name>OUT_0</name></connection>
<intersection>-121 9</intersection>
<intersection>-74.5 3</intersection>
<intersection>-63.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-63.5,72,-63.5</points>
<connection>
<GID>525</GID>
<name>IN_2</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>62.5,-74.5,72,-74.5</points>
<connection>
<GID>527</GID>
<name>IN_2</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>62.5,-121,72.5,-121</points>
<connection>
<GID>538</GID>
<name>IN_2</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-40.5,29,-40</points>
<intersection>-40.5 3</intersection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-40,33,-40</points>
<connection>
<GID>509</GID>
<name>IN_0</name></connection>
<intersection>27.5 4</intersection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>27.5,-40.5,29,-40.5</points>
<connection>
<GID>507</GID>
<name>OUT_0</name></connection>
<intersection>29 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>27.5,-129.5,27.5,-40</points>
<intersection>-129.5 15</intersection>
<intersection>-117 13</intersection>
<intersection>-105.5 11</intersection>
<intersection>-81 7</intersection>
<intersection>-70.5 5</intersection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>27.5,-70.5,72,-70.5</points>
<connection>
<GID>527</GID>
<name>IN_0</name></connection>
<intersection>27.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>27.5,-81,72,-81</points>
<connection>
<GID>529</GID>
<name>IN_0</name></connection>
<intersection>27.5 4</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>27.5,-105.5,72,-105.5</points>
<connection>
<GID>537</GID>
<name>IN_0</name></connection>
<intersection>27.5 4</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>27.5,-117,72.5,-117</points>
<connection>
<GID>538</GID>
<name>IN_0</name></connection>
<intersection>27.5 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>27.5,-129.5,72.5,-129.5</points>
<connection>
<GID>539</GID>
<name>IN_0</name></connection>
<intersection>27.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-58,84.5,-48</points>
<intersection>-58 2</intersection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,-48,84.5,-48</points>
<connection>
<GID>523</GID>
<name>OUT</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-58,91,-58</points>
<connection>
<GID>535</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-61.5,84.5,-60</points>
<intersection>-61.5 2</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84.5,-60,91,-60</points>
<connection>
<GID>535</GID>
<name>IN_1</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78,-61.5,84.5,-61.5</points>
<connection>
<GID>525</GID>
<name>OUT</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-72.5,84.5,-62</points>
<intersection>-72.5 2</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84.5,-62,91,-62</points>
<connection>
<GID>535</GID>
<name>IN_2</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78,-72.5,84.5,-72.5</points>
<connection>
<GID>527</GID>
<name>OUT</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-83,90,-64</points>
<intersection>-83 2</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-64,91,-64</points>
<connection>
<GID>535</GID>
<name>IN_3</name></connection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78,-83,90,-83</points>
<connection>
<GID>529</GID>
<name>OUT</name></connection>
<intersection>90 0</intersection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-61,102,-59</points>
<intersection>-61 2</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102,-59,106.5,-59</points>
<connection>
<GID>533</GID>
<name>N_in0</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>98,-61,102,-61</points>
<connection>
<GID>535</GID>
<name>OUT</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,-104,105,-102</points>
<intersection>-104 2</intersection>
<intersection>-102 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-102,109.5,-102</points>
<connection>
<GID>543</GID>
<name>N_in0</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>101,-104,105,-104</points>
<connection>
<GID>544</GID>
<name>OUT</name></connection>
<intersection>105 0</intersection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-101,85.5,-95</points>
<intersection>-101 2</intersection>
<intersection>-95 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-95,85.5,-95</points>
<connection>
<GID>536</GID>
<name>OUT</name></connection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85.5,-101,94,-101</points>
<connection>
<GID>544</GID>
<name>IN_0</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-107.5,86,-103</points>
<intersection>-107.5 1</intersection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,-107.5,86,-107.5</points>
<connection>
<GID>537</GID>
<name>OUT</name></connection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86,-103,94,-103</points>
<connection>
<GID>544</GID>
<name>IN_1</name></connection>
<intersection>86 0</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-119,86,-105</points>
<intersection>-119 1</intersection>
<intersection>-105 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78.5,-119,86,-119</points>
<connection>
<GID>538</GID>
<name>OUT</name></connection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86,-105,94,-105</points>
<connection>
<GID>544</GID>
<name>IN_2</name></connection>
<intersection>86 0</intersection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-131.5,86,-107</points>
<intersection>-131.5 1</intersection>
<intersection>-107 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78.5,-131.5,86,-131.5</points>
<connection>
<GID>539</GID>
<name>OUT</name></connection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86,-107,94,-107</points>
<connection>
<GID>544</GID>
<name>IN_3</name></connection>
<intersection>86 0</intersection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>